----------------------------------------------------------------------------------------------------
-- Copyright (c) 2019 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- This is a single-ported ROM (Wishbone B4 pipelined interface).
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
  port(
    -- Control signals.
    i_clk : in std_logic;

    -- Wishbone memory interface (b4 pipelined slave).
    -- See: https://cdn.opencores.org/downloads/wbspec_b4.pdf
    i_wb_cyc : in std_logic;
    i_wb_stb : in std_logic;
    i_wb_adr : in std_logic_vector(31 downto 2);
    o_wb_dat : out std_logic_vector(31 downto 0);
    o_wb_ack : out std_logic;
    o_wb_stall : out std_logic
  );
end rom;

architecture rtl of rom is
  constant C_ADDR_BITS : positive := 11;

  signal s_is_valid_wb_request : std_logic;
  signal s_rom_addr : std_logic_vector(C_ADDR_BITS-1 downto 0);
begin
  -- Wishbone control logic.
  s_is_valid_wb_request <= i_wb_cyc and i_wb_stb;

  -- We always ack and never stall - we're that fast ;-)
  process(i_clk)
  begin
    if rising_edge(i_clk) then
      o_wb_ack <= s_is_valid_wb_request;
    end if;
  end process;
  o_wb_stall <= '0';

  -- Actual ROM.
  s_rom_addr <= i_wb_adr(C_ADDR_BITS+1 downto 2);

  process(i_clk)
  begin
    if rising_edge(i_clk) then
      case s_rom_addr is
        when 11x"0" => o_wb_dat <= x"00000000";
        when 11x"1" => o_wb_dat <= x"00000000";
        when 11x"2" => o_wb_dat <= x"00000000";
        when 11x"3" => o_wb_dat <= x"00000000";
        when 11x"4" => o_wb_dat <= x"00000000";
        when 11x"5" => o_wb_dat <= x"00000000";
        when 11x"6" => o_wb_dat <= x"00000000";
        when 11x"7" => o_wb_dat <= x"00000000";
        when 11x"8" => o_wb_dat <= x"00000000";
        when 11x"9" => o_wb_dat <= x"00000000";
        when 11x"a" => o_wb_dat <= x"00000000";
        when 11x"b" => o_wb_dat <= x"00000000";
        when 11x"c" => o_wb_dat <= x"00000000";
        when 11x"d" => o_wb_dat <= x"00000000";
        when 11x"e" => o_wb_dat <= x"00000000";
        when 11x"f" => o_wb_dat <= x"00000000";
        when 11x"10" => o_wb_dat <= x"00000000";
        when 11x"11" => o_wb_dat <= x"00000000";
        when 11x"12" => o_wb_dat <= x"00000000";
        when 11x"13" => o_wb_dat <= x"00000000";
        when 11x"14" => o_wb_dat <= x"00000000";
        when 11x"15" => o_wb_dat <= x"00000000";
        when 11x"16" => o_wb_dat <= x"00000000";
        when 11x"17" => o_wb_dat <= x"00000000";
        when 11x"18" => o_wb_dat <= x"00000000";
        when 11x"19" => o_wb_dat <= x"00000000";
        when 11x"1a" => o_wb_dat <= x"00000000";
        when 11x"1b" => o_wb_dat <= x"00000000";
        when 11x"1c" => o_wb_dat <= x"00000000";
        when 11x"1d" => o_wb_dat <= x"00000000";
        when 11x"1e" => o_wb_dat <= x"00000000";
        when 11x"1f" => o_wb_dat <= x"00000000";
        when 11x"20" => o_wb_dat <= x"00000000";
        when 11x"21" => o_wb_dat <= x"00000000";
        when 11x"22" => o_wb_dat <= x"00000000";
        when 11x"23" => o_wb_dat <= x"00000000";
        when 11x"24" => o_wb_dat <= x"00000000";
        when 11x"25" => o_wb_dat <= x"00000000";
        when 11x"26" => o_wb_dat <= x"00000000";
        when 11x"27" => o_wb_dat <= x"00000000";
        when 11x"28" => o_wb_dat <= x"00000000";
        when 11x"29" => o_wb_dat <= x"00000000";
        when 11x"2a" => o_wb_dat <= x"00000000";
        when 11x"2b" => o_wb_dat <= x"00000000";
        when 11x"2c" => o_wb_dat <= x"00000000";
        when 11x"2d" => o_wb_dat <= x"00000000";
        when 11x"2e" => o_wb_dat <= x"00000000";
        when 11x"2f" => o_wb_dat <= x"00000000";
        when 11x"30" => o_wb_dat <= x"00000000";
        when 11x"31" => o_wb_dat <= x"00000000";
        when 11x"32" => o_wb_dat <= x"00000000";
        when 11x"33" => o_wb_dat <= x"00000000";
        when 11x"34" => o_wb_dat <= x"00000000";
        when 11x"35" => o_wb_dat <= x"00000000";
        when 11x"36" => o_wb_dat <= x"00000000";
        when 11x"37" => o_wb_dat <= x"00000000";
        when 11x"38" => o_wb_dat <= x"00000000";
        when 11x"39" => o_wb_dat <= x"00000000";
        when 11x"3a" => o_wb_dat <= x"00000000";
        when 11x"3b" => o_wb_dat <= x"00000000";
        when 11x"3c" => o_wb_dat <= x"00000000";
        when 11x"3d" => o_wb_dat <= x"00000000";
        when 11x"3e" => o_wb_dat <= x"00000000";
        when 11x"3f" => o_wb_dat <= x"00000000";
        when 11x"40" => o_wb_dat <= x"00000000";
        when 11x"41" => o_wb_dat <= x"00000000";
        when 11x"42" => o_wb_dat <= x"00000000";
        when 11x"43" => o_wb_dat <= x"00000000";
        when 11x"44" => o_wb_dat <= x"00000000";
        when 11x"45" => o_wb_dat <= x"00000000";
        when 11x"46" => o_wb_dat <= x"00000000";
        when 11x"47" => o_wb_dat <= x"00000000";
        when 11x"48" => o_wb_dat <= x"00000000";
        when 11x"49" => o_wb_dat <= x"00000000";
        when 11x"4a" => o_wb_dat <= x"00000000";
        when 11x"4b" => o_wb_dat <= x"00000000";
        when 11x"4c" => o_wb_dat <= x"00000000";
        when 11x"4d" => o_wb_dat <= x"00000000";
        when 11x"4e" => o_wb_dat <= x"00000000";
        when 11x"4f" => o_wb_dat <= x"00000000";
        when 11x"50" => o_wb_dat <= x"00000000";
        when 11x"51" => o_wb_dat <= x"00000000";
        when 11x"52" => o_wb_dat <= x"00000000";
        when 11x"53" => o_wb_dat <= x"00000000";
        when 11x"54" => o_wb_dat <= x"00000000";
        when 11x"55" => o_wb_dat <= x"00000000";
        when 11x"56" => o_wb_dat <= x"00000000";
        when 11x"57" => o_wb_dat <= x"00000000";
        when 11x"58" => o_wb_dat <= x"00000000";
        when 11x"59" => o_wb_dat <= x"00000000";
        when 11x"5a" => o_wb_dat <= x"00000000";
        when 11x"5b" => o_wb_dat <= x"00000000";
        when 11x"5c" => o_wb_dat <= x"00000000";
        when 11x"5d" => o_wb_dat <= x"00000000";
        when 11x"5e" => o_wb_dat <= x"00000000";
        when 11x"5f" => o_wb_dat <= x"00000000";
        when 11x"60" => o_wb_dat <= x"00000000";
        when 11x"61" => o_wb_dat <= x"00000000";
        when 11x"62" => o_wb_dat <= x"00000000";
        when 11x"63" => o_wb_dat <= x"00000000";
        when 11x"64" => o_wb_dat <= x"00000000";
        when 11x"65" => o_wb_dat <= x"00000000";
        when 11x"66" => o_wb_dat <= x"00000000";
        when 11x"67" => o_wb_dat <= x"00000000";
        when 11x"68" => o_wb_dat <= x"00000000";
        when 11x"69" => o_wb_dat <= x"00000000";
        when 11x"6a" => o_wb_dat <= x"00000000";
        when 11x"6b" => o_wb_dat <= x"00000000";
        when 11x"6c" => o_wb_dat <= x"00000000";
        when 11x"6d" => o_wb_dat <= x"00000000";
        when 11x"6e" => o_wb_dat <= x"00000000";
        when 11x"6f" => o_wb_dat <= x"00000000";
        when 11x"70" => o_wb_dat <= x"00000000";
        when 11x"71" => o_wb_dat <= x"00000000";
        when 11x"72" => o_wb_dat <= x"00000000";
        when 11x"73" => o_wb_dat <= x"00000000";
        when 11x"74" => o_wb_dat <= x"00000000";
        when 11x"75" => o_wb_dat <= x"00000000";
        when 11x"76" => o_wb_dat <= x"00000000";
        when 11x"77" => o_wb_dat <= x"00000000";
        when 11x"78" => o_wb_dat <= x"00000000";
        when 11x"79" => o_wb_dat <= x"00000000";
        when 11x"7a" => o_wb_dat <= x"00000000";
        when 11x"7b" => o_wb_dat <= x"00000000";
        when 11x"7c" => o_wb_dat <= x"00000000";
        when 11x"7d" => o_wb_dat <= x"00000000";
        when 11x"7e" => o_wb_dat <= x"00000000";
        when 11x"7f" => o_wb_dat <= x"00000000";
        when 11x"80" => o_wb_dat <= x"ec400000";
        when 11x"81" => o_wb_dat <= x"40420078";
        when 11x"82" => o_wb_dat <= x"c040000a";
        when 11x"83" => o_wb_dat <= x"8c420002";
        when 11x"84" => o_wb_dat <= x"ec280000";
        when 11x"85" => o_wb_dat <= x"40210100";
        when 11x"86" => o_wb_dat <= x"00600000";
        when 11x"87" => o_wb_dat <= x"03a2061d";
        when 11x"88" => o_wb_dat <= x"2c018004";
        when 11x"89" => o_wb_dat <= x"005d0416";
        when 11x"8a" => o_wb_dat <= x"00213b07";
        when 11x"8b" => o_wb_dat <= x"c45ffffc";
        when 11x"8c" => o_wb_dat <= x"ec380000";
        when 11x"8d" => o_wb_dat <= x"0c21000c";
        when 11x"8e" => o_wb_dat <= x"ef880000";
        when 11x"8f" => o_wb_dat <= x"039c0215";
        when 11x"90" => o_wb_dat <= x"e7e00269";
        when 11x"91" => o_wb_dat <= x"02a00210";
        when 11x"92" => o_wb_dat <= x"ec580000";
        when 11x"93" => o_wb_dat <= x"0c42000c";
        when 11x"94" => o_wb_dat <= x"ec680000";
        when 11x"95" => o_wb_dat <= x"00630415";
        when 11x"96" => o_wb_dat <= x"e8401000";
        when 11x"97" => o_wb_dat <= x"00410415";
        when 11x"98" => o_wb_dat <= x"02820616";
        when 11x"99" => o_wb_dat <= x"00202810";
        when 11x"9a" => o_wb_dat <= x"e7e00261";
        when 11x"9b" => o_wb_dat <= x"1c3f14f4";
        when 11x"9c" => o_wb_dat <= x"e7e002b1";
        when 11x"9d" => o_wb_dat <= x"1c3f1509";
        when 11x"9e" => o_wb_dat <= x"ec480000";
        when 11x"9f" => o_wb_dat <= x"ec780000";
        when 11x"a0" => o_wb_dat <= x"0c63000c";
        when 11x"a1" => o_wb_dat <= x"e7e0006f";
        when 11x"a2" => o_wb_dat <= x"1c3f14ff";
        when 11x"a3" => o_wb_dat <= x"ec500000";
        when 11x"a4" => o_wb_dat <= x"ec780000";
        when 11x"a5" => o_wb_dat <= x"0c630010";
        when 11x"a6" => o_wb_dat <= x"e7e0006a";
        when 11x"a7" => o_wb_dat <= x"1c3f14f5";
        when 11x"a8" => o_wb_dat <= x"ec480000";
        when 11x"a9" => o_wb_dat <= x"40420100";
        when 11x"aa" => o_wb_dat <= x"ec600000";
        when 11x"ab" => o_wb_dat <= x"40630078";
        when 11x"ac" => o_wb_dat <= x"e7e00064";
        when 11x"ad" => o_wb_dat <= x"1c3f14e7";
        when 11x"ae" => o_wb_dat <= x"00402810";
        when 11x"af" => o_wb_dat <= x"00602a10";
        when 11x"b0" => o_wb_dat <= x"e7e00060";
        when 11x"b1" => o_wb_dat <= x"1c3f14e1";
        when 11x"b2" => o_wb_dat <= x"e8601000";
        when 11x"b3" => o_wb_dat <= x"00403810";
        when 11x"b4" => o_wb_dat <= x"00430416";
        when 11x"b5" => o_wb_dat <= x"e7e0005b";
        when 11x"b6" => o_wb_dat <= x"e7e00177";
        when 11x"b7" => o_wb_dat <= x"ec300000";
        when 11x"b8" => o_wb_dat <= x"40210000";
        when 11x"b9" => o_wb_dat <= x"ec580000";
        when 11x"ba" => o_wb_dat <= x"0c420010";
        when 11x"bb" => o_wb_dat <= x"e8600002";
        when 11x"bc" => o_wb_dat <= x"e7e00174";
        when 11x"bd" => o_wb_dat <= x"ec280000";
        when 11x"be" => o_wb_dat <= x"40210178";
        when 11x"bf" => o_wb_dat <= x"00412816";
        when 11x"c0" => o_wb_dat <= x"e8600001";
        when 11x"c1" => o_wb_dat <= x"e7e0016f";
        when 11x"c2" => o_wb_dat <= x"1c3f14b2";
        when 11x"c3" => o_wb_dat <= x"e7e0028a";
        when 11x"c4" => o_wb_dat <= x"e8200000";
        when 11x"c5" => o_wb_dat <= x"e8400000";
        when 11x"c6" => o_wb_dat <= x"e8600000";
        when 11x"c7" => o_wb_dat <= x"e8800000";
        when 11x"c8" => o_wb_dat <= x"e8a00000";
        when 11x"c9" => o_wb_dat <= x"e8c00000";
        when 11x"ca" => o_wb_dat <= x"e8e00000";
        when 11x"cb" => o_wb_dat <= x"e9000000";
        when 11x"cc" => o_wb_dat <= x"e9200000";
        when 11x"cd" => o_wb_dat <= x"e9400000";
        when 11x"ce" => o_wb_dat <= x"e9600000";
        when 11x"cf" => o_wb_dat <= x"e9800000";
        when 11x"d0" => o_wb_dat <= x"e9a00000";
        when 11x"d1" => o_wb_dat <= x"e9c00000";
        when 11x"d2" => o_wb_dat <= x"e9e00000";
        when 11x"d3" => o_wb_dat <= x"ea000000";
        when 11x"d4" => o_wb_dat <= x"ea200000";
        when 11x"d5" => o_wb_dat <= x"ea400000";
        when 11x"d6" => o_wb_dat <= x"ea600000";
        when 11x"d7" => o_wb_dat <= x"ea800000";
        when 11x"d8" => o_wb_dat <= x"eaa00000";
        when 11x"d9" => o_wb_dat <= x"eac00000";
        when 11x"da" => o_wb_dat <= x"eae00000";
        when 11x"db" => o_wb_dat <= x"eb000000";
        when 11x"dc" => o_wb_dat <= x"eb200000";
        when 11x"dd" => o_wb_dat <= x"eb400000";
        when 11x"de" => o_wb_dat <= x"eb600000";
        when 11x"df" => o_wb_dat <= x"eba00000";
        when 11x"e0" => o_wb_dat <= x"ebc00000";
        when 11x"e1" => o_wb_dat <= x"03a00000";
        when 11x"e2" => o_wb_dat <= x"40208000";
        when 11x"e3" => o_wb_dat <= x"40408000";
        when 11x"e4" => o_wb_dat <= x"40608000";
        when 11x"e5" => o_wb_dat <= x"40808000";
        when 11x"e6" => o_wb_dat <= x"40a08000";
        when 11x"e7" => o_wb_dat <= x"40c08000";
        when 11x"e8" => o_wb_dat <= x"40e08000";
        when 11x"e9" => o_wb_dat <= x"41008000";
        when 11x"ea" => o_wb_dat <= x"41208000";
        when 11x"eb" => o_wb_dat <= x"41408000";
        when 11x"ec" => o_wb_dat <= x"41608000";
        when 11x"ed" => o_wb_dat <= x"41808000";
        when 11x"ee" => o_wb_dat <= x"41a08000";
        when 11x"ef" => o_wb_dat <= x"41c08000";
        when 11x"f0" => o_wb_dat <= x"41e08000";
        when 11x"f1" => o_wb_dat <= x"42008000";
        when 11x"f2" => o_wb_dat <= x"42208000";
        when 11x"f3" => o_wb_dat <= x"42408000";
        when 11x"f4" => o_wb_dat <= x"42608000";
        when 11x"f5" => o_wb_dat <= x"42808000";
        when 11x"f6" => o_wb_dat <= x"42a08000";
        when 11x"f7" => o_wb_dat <= x"42c08000";
        when 11x"f8" => o_wb_dat <= x"42e08000";
        when 11x"f9" => o_wb_dat <= x"43008000";
        when 11x"fa" => o_wb_dat <= x"43208000";
        when 11x"fb" => o_wb_dat <= x"43408000";
        when 11x"fc" => o_wb_dat <= x"43608000";
        when 11x"fd" => o_wb_dat <= x"43808000";
        when 11x"fe" => o_wb_dat <= x"43a08000";
        when 11x"ff" => o_wb_dat <= x"43c08000";
        when 11x"100" => o_wb_dat <= x"43e08000";
        when 11x"101" => o_wb_dat <= x"e8200001";
        when 11x"102" => o_wb_dat <= x"ec400002";
        when 11x"103" => o_wb_dat <= x"54420754";
        when 11x"104" => o_wb_dat <= x"e7e00020";
        when 11x"105" => o_wb_dat <= x"00000000";
        when 11x"106" => o_wb_dat <= x"00000000";
        when 11x"107" => o_wb_dat <= x"00000000";
        when 11x"108" => o_wb_dat <= x"00000000";
        when 11x"109" => o_wb_dat <= x"00000000";
        when 11x"10a" => o_wb_dat <= x"e3e00000";
        when 11x"10b" => o_wb_dat <= x"00000000";
        when 11x"10c" => o_wb_dat <= x"00000000";
        when 11x"10d" => o_wb_dat <= x"00000000";
        when 11x"10e" => o_wb_dat <= x"00000000";
        when 11x"10f" => o_wb_dat <= x"00000000";
        when 11x"110" => o_wb_dat <= x"579c7ff4";
        when 11x"111" => o_wb_dat <= x"2fdc0000";
        when 11x"112" => o_wb_dat <= x"2e9c0004";
        when 11x"113" => o_wb_dat <= x"2ebc0008";
        when 11x"114" => o_wb_dat <= x"02800410";
        when 11x"115" => o_wb_dat <= x"02a00610";
        when 11x"116" => o_wb_dat <= x"e7e00237";
        when 11x"117" => o_wb_dat <= x"00202810";
        when 11x"118" => o_wb_dat <= x"e7e00279";
        when 11x"119" => o_wb_dat <= x"1c3f134b";
        when 11x"11a" => o_wb_dat <= x"e7e00233";
        when 11x"11b" => o_wb_dat <= x"00202a10";
        when 11x"11c" => o_wb_dat <= x"e7e00286";
        when 11x"11d" => o_wb_dat <= x"1c3f133e";
        when 11x"11e" => o_wb_dat <= x"e7e0022f";
        when 11x"11f" => o_wb_dat <= x"0fdc0000";
        when 11x"120" => o_wb_dat <= x"0e9c0004";
        when 11x"121" => o_wb_dat <= x"0ebc0008";
        when 11x"122" => o_wb_dat <= x"579c000c";
        when 11x"123" => o_wb_dat <= x"e3c00000";
        when 11x"124" => o_wb_dat <= x"579c7ffc";
        when 11x"125" => o_wb_dat <= x"2fdc0000";
        when 11x"126" => o_wb_dat <= x"e7e00005";
        when 11x"127" => o_wb_dat <= x"e7e0005e";
        when 11x"128" => o_wb_dat <= x"0fdc0000";
        when 11x"129" => o_wb_dat <= x"579c0004";
        when 11x"12a" => o_wb_dat <= x"e3c00000";
        when 11x"12b" => o_wb_dat <= x"579c7ffc";
        when 11x"12c" => o_wb_dat <= x"2fbc0000";
        when 11x"12d" => o_wb_dat <= x"ed680000";
        when 11x"12e" => o_wb_dat <= x"416b0000";
        when 11x"12f" => o_wb_dat <= x"ed90400a";
        when 11x"130" => o_wb_dat <= x"418c0555";
        when 11x"131" => o_wb_dat <= x"2d8b0000";
        when 11x"132" => o_wb_dat <= x"ed90a000";
        when 11x"133" => o_wb_dat <= x"418c0002";
        when 11x"134" => o_wb_dat <= x"2d8b0004";
        when 11x"135" => o_wb_dat <= x"ed90c000";
        when 11x"136" => o_wb_dat <= x"418c0001";
        when 11x"137" => o_wb_dat <= x"2d8b0008";
        when 11x"138" => o_wb_dat <= x"ed8c0000";
        when 11x"139" => o_wb_dat <= x"418c00ff";
        when 11x"13a" => o_wb_dat <= x"2d8b000c";
        when 11x"13b" => o_wb_dat <= x"556b0010";
        when 11x"13c" => o_wb_dat <= x"e8200064";
        when 11x"13d" => o_wb_dat <= x"e8400032";
        when 11x"13e" => o_wb_dat <= x"e8600000";
        when 11x"13f" => o_wb_dat <= x"e8800002";
        when 11x"140" => o_wb_dat <= x"e8a00003";
        when 11x"141" => o_wb_dat <= x"e8c00001";
        when 11x"142" => o_wb_dat <= x"edffe000";
        when 11x"143" => o_wb_dat <= x"2deb0000";
        when 11x"144" => o_wb_dat <= x"e9c00001";
        when 11x"145" => o_wb_dat <= x"88e30010";
        when 11x"146" => o_wb_dat <= x"89020008";
        when 11x"147" => o_wb_dat <= x"00e71010";
        when 11x"148" => o_wb_dat <= x"00e70210";
        when 11x"149" => o_wb_dat <= x"00e71e10";
        when 11x"14a" => o_wb_dat <= x"00eb1d0b";
        when 11x"14b" => o_wb_dat <= x"00210815";
        when 11x"14c" => o_wb_dat <= x"6ce100ff";
        when 11x"14d" => o_wb_dat <= x"0100021b";
        when 11x"14e" => o_wb_dat <= x"00e71012";
        when 11x"14f" => o_wb_dat <= x"c8e00003";
        when 11x"150" => o_wb_dat <= x"00840016";
        when 11x"151" => o_wb_dat <= x"00210815";
        when 11x"152" => o_wb_dat <= x"00420a15";
        when 11x"153" => o_wb_dat <= x"6ce200ff";
        when 11x"154" => o_wb_dat <= x"0100041b";
        when 11x"155" => o_wb_dat <= x"00e71012";
        when 11x"156" => o_wb_dat <= x"c8e00003";
        when 11x"157" => o_wb_dat <= x"00a50016";
        when 11x"158" => o_wb_dat <= x"00420a15";
        when 11x"159" => o_wb_dat <= x"00630c15";
        when 11x"15a" => o_wb_dat <= x"6ce300ff";
        when 11x"15b" => o_wb_dat <= x"0100061b";
        when 11x"15c" => o_wb_dat <= x"00e71012";
        when 11x"15d" => o_wb_dat <= x"c8e00003";
        when 11x"15e" => o_wb_dat <= x"00c60016";
        when 11x"15f" => o_wb_dat <= x"00630c15";
        when 11x"160" => o_wb_dat <= x"55ce0001";
        when 11x"161" => o_wb_dat <= x"60ee0100";
        when 11x"162" => o_wb_dat <= x"c8ffffe3";
        when 11x"163" => o_wb_dat <= x"556b0400";
        when 11x"164" => o_wb_dat <= x"ec2a0000";
        when 11x"165" => o_wb_dat <= x"ec500000";
        when 11x"166" => o_wb_dat <= x"40420400";
        when 11x"167" => o_wb_dat <= x"2c2b0000";
        when 11x"168" => o_wb_dat <= x"2c4b0004";
        when 11x"169" => o_wb_dat <= x"ed908000";
        when 11x"16a" => o_wb_dat <= x"418c0780";
        when 11x"16b" => o_wb_dat <= x"2d8b0008";
        when 11x"16c" => o_wb_dat <= x"556b000c";
        when 11x"16d" => o_wb_dat <= x"e3e00004";
        when 11x"16e" => o_wb_dat <= x"2c2b0000";
        when 11x"16f" => o_wb_dat <= x"2c4b0004";
        when 11x"170" => o_wb_dat <= x"556b0008";
        when 11x"171" => o_wb_dat <= x"54210003";
        when 11x"172" => o_wb_dat <= x"544200a0";
        when 11x"173" => o_wb_dat <= x"49a13fff";
        when 11x"174" => o_wb_dat <= x"65ad0438";
        when 11x"175" => o_wb_dat <= x"c9bffff9";
        when 11x"176" => o_wb_dat <= x"ed8a000f";
        when 11x"177" => o_wb_dat <= x"418c07ff";
        when 11x"178" => o_wb_dat <= x"2d8b0000";
        when 11x"179" => o_wb_dat <= x"ed280002";
        when 11x"17a" => o_wb_dat <= x"41290000";
        when 11x"17b" => o_wb_dat <= x"01400000";
        when 11x"17c" => o_wb_dat <= x"e960e100";
        when 11x"17d" => o_wb_dat <= x"03aa161d";
        when 11x"17e" => o_wb_dat <= x"017d1616";
        when 11x"17f" => o_wb_dat <= x"2c098004";
        when 11x"180" => o_wb_dat <= x"01293b07";
        when 11x"181" => o_wb_dat <= x"c57ffffc";
        when 11x"182" => o_wb_dat <= x"0fbc0000";
        when 11x"183" => o_wb_dat <= x"579c0004";
        when 11x"184" => o_wb_dat <= x"e3c00000";
        when 11x"185" => o_wb_dat <= x"579c7ff4";
        when 11x"186" => o_wb_dat <= x"2fdc0000";
        when 11x"187" => o_wb_dat <= x"2e9c0004";
        when 11x"188" => o_wb_dat <= x"2ebc0008";
        when 11x"189" => o_wb_dat <= x"ee980000";
        when 11x"18a" => o_wb_dat <= x"eaa00001";
        when 11x"18b" => o_wb_dat <= x"00202a10";
        when 11x"18c" => o_wb_dat <= x"e7e0000f";
        when 11x"18d" => o_wb_dat <= x"0c340024";
        when 11x"18e" => o_wb_dat <= x"e7e00086";
        when 11x"18f" => o_wb_dat <= x"2eb40060";
        when 11x"190" => o_wb_dat <= x"0c540020";
        when 11x"191" => o_wb_dat <= x"0c340020";
        when 11x"192" => o_wb_dat <= x"00210418";
        when 11x"193" => o_wb_dat <= x"cc3ffffe";
        when 11x"194" => o_wb_dat <= x"56b50001";
        when 11x"195" => o_wb_dat <= x"e3fffff6";
        when 11x"196" => o_wb_dat <= x"0fdc0000";
        when 11x"197" => o_wb_dat <= x"0e9c0004";
        when 11x"198" => o_wb_dat <= x"0ebc0008";
        when 11x"199" => o_wb_dat <= x"579c000c";
        when 11x"19a" => o_wb_dat <= x"e3c00000";
        when 11x"19b" => o_wb_dat <= x"579c7ffc";
        when 11x"19c" => o_wb_dat <= x"2fdc0000";
        when 11x"19d" => o_wb_dat <= x"ec580000";
        when 11x"19e" => o_wb_dat <= x"0c420028";
        when 11x"19f" => o_wb_dat <= x"48420001";
        when 11x"1a0" => o_wb_dat <= x"c0400003";
        when 11x"1a1" => o_wb_dat <= x"e7e00043";
        when 11x"1a2" => o_wb_dat <= x"c0000002";
        when 11x"1a3" => o_wb_dat <= x"e7e00004";
        when 11x"1a4" => o_wb_dat <= x"0fdc0000";
        when 11x"1a5" => o_wb_dat <= x"579c0004";
        when 11x"1a6" => o_wb_dat <= x"e3c00000";
        when 11x"1a7" => o_wb_dat <= x"579c7ffc";
        when 11x"1a8" => o_wb_dat <= x"2e9c0000";
        when 11x"1a9" => o_wb_dat <= x"0dbf00e8";
        when 11x"1aa" => o_wb_dat <= x"0e3f00d4";
        when 11x"1ab" => o_wb_dat <= x"0e5f00d4";
        when 11x"1ac" => o_wb_dat <= x"00210068";
        when 11x"1ad" => o_wb_dat <= x"00210272";
        when 11x"1ae" => o_wb_dat <= x"ec478478";
        when 11x"1af" => o_wb_dat <= x"00410472";
        when 11x"1b0" => o_wb_dat <= x"ec67f000";
        when 11x"1b1" => o_wb_dat <= x"00420670";
        when 11x"1b2" => o_wb_dat <= x"02830473";
        when 11x"1b3" => o_wb_dat <= x"01ad2872";
        when 11x"1b4" => o_wb_dat <= x"edc80002";
        when 11x"1b5" => o_wb_dat <= x"41ce0000";
        when 11x"1b6" => o_wb_dat <= x"ea000168";
        when 11x"1b7" => o_wb_dat <= x"84700001";
        when 11x"1b8" => o_wb_dat <= x"00630068";
        when 11x"1b9" => o_wb_dat <= x"006d0672";
        when 11x"1ba" => o_wb_dat <= x"0c5f00a0";
        when 11x"1bb" => o_wb_dat <= x"00420671";
        when 11x"1bc" => o_wb_dat <= x"e9e00280";
        when 11x"1bd" => o_wb_dat <= x"846f0001";
        when 11x"1be" => o_wb_dat <= x"00630068";
        when 11x"1bf" => o_wb_dat <= x"006d0672";
        when 11x"1c0" => o_wb_dat <= x"0c3f0084";
        when 11x"1c1" => o_wb_dat <= x"00210671";
        when 11x"1c2" => o_wb_dat <= x"00600010";
        when 11x"1c3" => o_wb_dat <= x"00800010";
        when 11x"1c4" => o_wb_dat <= x"e9200000";
        when 11x"1c5" => o_wb_dat <= x"00a30672";
        when 11x"1c6" => o_wb_dat <= x"00c40872";
        when 11x"1c7" => o_wb_dat <= x"55290001";
        when 11x"1c8" => o_wb_dat <= x"00830872";
        when 11x"1c9" => o_wb_dat <= x"00650c71";
        when 11x"1ca" => o_wb_dat <= x"00a50c70";
        when 11x"1cb" => o_wb_dat <= x"00840870";
        when 11x"1cc" => o_wb_dat <= x"00630270";
        when 11x"1cd" => o_wb_dat <= x"01492219";
        when 11x"1ce" => o_wb_dat <= x"00840470";
        when 11x"1cf" => o_wb_dat <= x"00a52464";
        when 11x"1d0" => o_wb_dat <= x"cca00003";
        when 11x"1d1" => o_wb_dat <= x"c95ffff4";
        when 11x"1d2" => o_wb_dat <= x"e9200000";
        when 11x"1d3" => o_wb_dat <= x"89290001";
        when 11x"1d4" => o_wb_dat <= x"252e0000";
        when 11x"1d5" => o_wb_dat <= x"55ce0001";
        when 11x"1d6" => o_wb_dat <= x"55ef7fff";
        when 11x"1d7" => o_wb_dat <= x"00211a70";
        when 11x"1d8" => o_wb_dat <= x"ddffffea";
        when 11x"1d9" => o_wb_dat <= x"56107fff";
        when 11x"1da" => o_wb_dat <= x"00421a70";
        when 11x"1db" => o_wb_dat <= x"de1fffe1";
        when 11x"1dc" => o_wb_dat <= x"0e9c0000";
        when 11x"1dd" => o_wb_dat <= x"579c0004";
        when 11x"1de" => o_wb_dat <= x"e3c00000";
        when 11x"1df" => o_wb_dat <= x"0000007f";
        when 11x"1e0" => o_wb_dat <= x"40800000";
        when 11x"1e1" => o_wb_dat <= x"bf9403b1";
        when 11x"1e2" => o_wb_dat <= x"be8ef344";
        when 11x"1e3" => o_wb_dat <= x"3be56042";
        when 11x"1e4" => o_wb_dat <= x"579c7ff8";
        when 11x"1e5" => o_wb_dat <= x"2e9c0000";
        when 11x"1e6" => o_wb_dat <= x"2ebc0004";
        when 11x"1e7" => o_wb_dat <= x"00210215";
        when 11x"1e8" => o_wb_dat <= x"01a00000";
        when 11x"1e9" => o_wb_dat <= x"03a01a10";
        when 11x"1ea" => o_wb_dat <= x"544d7fff";
        when 11x"1eb" => o_wb_dat <= x"1c82ffff";
        when 11x"1ec" => o_wb_dat <= x"eea00001";
        when 11x"1ed" => o_wb_dat <= x"42b50754";
        when 11x"1ee" => o_wb_dat <= x"ecc80002";
        when 11x"1ef" => o_wb_dat <= x"40c60000";
        when 11x"1f0" => o_wb_dat <= x"e9000168";
        when 11x"1f1" => o_wb_dat <= x"55087fff";
        when 11x"1f2" => o_wb_dat <= x"01280215";
        when 11x"1f3" => o_wb_dat <= x"e8e00140";
        when 11x"1f4" => o_wb_dat <= x"03ad0e1d";
        when 11x"1f5" => o_wb_dat <= x"00fd0e16";
        when 11x"1f6" => o_wb_dat <= x"00e48e15";
        when 11x"1f7" => o_wb_dat <= x"02870287";
        when 11x"1f8" => o_wb_dat <= x"0124a815";
        when 11x"1f9" => o_wb_dat <= x"490983ff";
        when 11x"1fa" => o_wb_dat <= x"0115d082";
        when 11x"1fb" => o_wb_dat <= x"00e7d140";
        when 11x"1fc" => o_wb_dat <= x"00279315";
        when 11x"1fd" => o_wb_dat <= x"2c268002";
        when 11x"1fe" => o_wb_dat <= x"00c61a87";
        when 11x"1ff" => o_wb_dat <= x"dcfffff5";
        when 11x"200" => o_wb_dat <= x"dd1ffff1";
        when 11x"201" => o_wb_dat <= x"0e9c0000";
        when 11x"202" => o_wb_dat <= x"0ebc0004";
        when 11x"203" => o_wb_dat <= x"579c0008";
        when 11x"204" => o_wb_dat <= x"e3c00000";
        when 11x"205" => o_wb_dat <= x"ec580000";
        when 11x"206" => o_wb_dat <= x"2c220060";
        when 11x"207" => o_wb_dat <= x"e3c00000";
        when 11x"208" => o_wb_dat <= x"1c5f0084";
        when 11x"209" => o_wb_dat <= x"ec780000";
        when 11x"20a" => o_wb_dat <= x"1c630040";
        when 11x"20b" => o_wb_dat <= x"e8a00008";
        when 11x"20c" => o_wb_dat <= x"4881000f";
        when 11x"20d" => o_wb_dat <= x"8c210004";
        when 11x"20e" => o_wb_dat <= x"00820805";
        when 11x"20f" => o_wb_dat <= x"2c830000";
        when 11x"210" => o_wb_dat <= x"54630004";
        when 11x"211" => o_wb_dat <= x"54a57fff";
        when 11x"212" => o_wb_dat <= x"c4bffffa";
        when 11x"213" => o_wb_dat <= x"e3c00000";
        when 11x"214" => o_wb_dat <= x"1c5f0054";
        when 11x"215" => o_wb_dat <= x"ec780000";
        when 11x"216" => o_wb_dat <= x"1c630040";
        when 11x"217" => o_wb_dat <= x"00e10019";
        when 11x"218" => o_wb_dat <= x"cce00003";
        when 11x"219" => o_wb_dat <= x"00210016";
        when 11x"21a" => o_wb_dat <= x"e8e00040";
        when 11x"21b" => o_wb_dat <= x"e8c0000a";
        when 11x"21c" => o_wb_dat <= x"e8a00008";
        when 11x"21d" => o_wb_dat <= x"00810c47";
        when 11x"21e" => o_wb_dat <= x"00210c45";
        when 11x"21f" => o_wb_dat <= x"00820805";
        when 11x"220" => o_wb_dat <= x"2c830000";
        when 11x"221" => o_wb_dat <= x"54630004";
        when 11x"222" => o_wb_dat <= x"54a57fff";
        when 11x"223" => o_wb_dat <= x"c0a00005";
        when 11x"224" => o_wb_dat <= x"c43ffff9";
        when 11x"225" => o_wb_dat <= x"00800e10";
        when 11x"226" => o_wb_dat <= x"e8e00000";
        when 11x"227" => o_wb_dat <= x"e3fffff9";
        when 11x"228" => o_wb_dat <= x"e3c00000";
        when 11x"229" => o_wb_dat <= x"4f5b063f";
        when 11x"22a" => o_wb_dat <= x"077d6d66";
        when 11x"22b" => o_wb_dat <= x"7c776f7f";
        when 11x"22c" => o_wb_dat <= x"71795e39";
        when 11x"22d" => o_wb_dat <= x"e8200000";
        when 11x"22e" => o_wb_dat <= x"2c3f7848";
        when 11x"22f" => o_wb_dat <= x"e3c00000";
        when 11x"230" => o_wb_dat <= x"0cbf7840";
        when 11x"231" => o_wb_dat <= x"6c850003";
        when 11x"232" => o_wb_dat <= x"cc800040";
        when 11x"233" => o_wb_dat <= x"8c820008";
        when 11x"234" => o_wb_dat <= x"78840080";
        when 11x"235" => o_wb_dat <= x"88c40004";
        when 11x"236" => o_wb_dat <= x"00c20c1a";
        when 11x"237" => o_wb_dat <= x"c8c0003b";
        when 11x"238" => o_wb_dat <= x"579c7fe8";
        when 11x"239" => o_wb_dat <= x"2e1c0014";
        when 11x"23a" => o_wb_dat <= x"2e3c0010";
        when 11x"23b" => o_wb_dat <= x"2e5c000c";
        when 11x"23c" => o_wb_dat <= x"2e7c0008";
        when 11x"23d" => o_wb_dat <= x"2e9c0004";
        when 11x"23e" => o_wb_dat <= x"2fdc0000";
        when 11x"23f" => o_wb_dat <= x"88c40003";
        when 11x"240" => o_wb_dat <= x"02050a15";
        when 11x"241" => o_wb_dat <= x"02100a15";
        when 11x"242" => o_wb_dat <= x"f4a7fffe";
        when 11x"243" => o_wb_dat <= x"54a507fc";
        when 11x"244" => o_wb_dat <= x"02052187";
        when 11x"245" => o_wb_dat <= x"2c900008";
        when 11x"246" => o_wb_dat <= x"e8800000";
        when 11x"247" => o_wb_dat <= x"2c90000c";
        when 11x"248" => o_wb_dat <= x"2c300014";
        when 11x"249" => o_wb_dat <= x"00210c15";
        when 11x"24a" => o_wb_dat <= x"2c300000";
        when 11x"24b" => o_wb_dat <= x"56900004";
        when 11x"24c" => o_wb_dat <= x"00460416";
        when 11x"24d" => o_wb_dat <= x"2c540000";
        when 11x"24e" => o_wb_dat <= x"56700010";
        when 11x"24f" => o_wb_dat <= x"2c730000";
        when 11x"250" => o_wb_dat <= x"f6200000";
        when 11x"251" => o_wb_dat <= x"563103f4";
        when 11x"252" => o_wb_dat <= x"f4200001";
        when 11x"253" => o_wb_dat <= x"542106d8";
        when 11x"254" => o_wb_dat <= x"e6200000";
        when 11x"255" => o_wb_dat <= x"f6400000";
        when 11x"256" => o_wb_dat <= x"565204f0";
        when 11x"257" => o_wb_dat <= x"0c300000";
        when 11x"258" => o_wb_dat <= x"e6400000";
        when 11x"259" => o_wb_dat <= x"f4200001";
        when 11x"25a" => o_wb_dat <= x"542106d0";
        when 11x"25b" => o_wb_dat <= x"e6200000";
        when 11x"25c" => o_wb_dat <= x"0c340000";
        when 11x"25d" => o_wb_dat <= x"f7c00000";
        when 11x"25e" => o_wb_dat <= x"e7c00145";
        when 11x"25f" => o_wb_dat <= x"f4200001";
        when 11x"260" => o_wb_dat <= x"542106bc";
        when 11x"261" => o_wb_dat <= x"e6200000";
        when 11x"262" => o_wb_dat <= x"0c330000";
        when 11x"263" => o_wb_dat <= x"e6400000";
        when 11x"264" => o_wb_dat <= x"f4200001";
        when 11x"265" => o_wb_dat <= x"542106c0";
        when 11x"266" => o_wb_dat <= x"e6200000";
        when 11x"267" => o_wb_dat <= x"0c3f7764";
        when 11x"268" => o_wb_dat <= x"54210001";
        when 11x"269" => o_wb_dat <= x"2c3f775c";
        when 11x"26a" => o_wb_dat <= x"0e1c0014";
        when 11x"26b" => o_wb_dat <= x"0e3c0010";
        when 11x"26c" => o_wb_dat <= x"0e5c000c";
        when 11x"26d" => o_wb_dat <= x"0e7c0008";
        when 11x"26e" => o_wb_dat <= x"0e9c0004";
        when 11x"26f" => o_wb_dat <= x"0fdc0000";
        when 11x"270" => o_wb_dat <= x"579c0018";
        when 11x"271" => o_wb_dat <= x"e3c00000";
        when 11x"272" => o_wb_dat <= x"e3c00000";
        when 11x"273" => o_wb_dat <= x"579c7ff8";
        when 11x"274" => o_wb_dat <= x"2e1c0004";
        when 11x"275" => o_wb_dat <= x"2fdc0000";
        when 11x"276" => o_wb_dat <= x"00600210";
        when 11x"277" => o_wb_dat <= x"f487fffe";
        when 11x"278" => o_wb_dat <= x"54840728";
        when 11x"279" => o_wb_dat <= x"e9800000";
        when 11x"27a" => o_wb_dat <= x"55610003";
        when 11x"27b" => o_wb_dat <= x"496b7ffc";
        when 11x"27c" => o_wb_dat <= x"e9bfffff";
        when 11x"27d" => o_wb_dat <= x"0c3f770c";
        when 11x"27e" => o_wb_dat <= x"002c021b";
        when 11x"27f" => o_wb_dat <= x"c8200003";
        when 11x"280" => o_wb_dat <= x"ea000000";
        when 11x"281" => o_wb_dat <= x"e3e00024";
        when 11x"282" => o_wb_dat <= x"0ca40010";
        when 11x"283" => o_wb_dat <= x"00220a12";
        when 11x"284" => o_wb_dat <= x"c020004b";
        when 11x"285" => o_wb_dat <= x"c060004a";
        when 11x"286" => o_wb_dat <= x"0cc4000c";
        when 11x"287" => o_wb_dat <= x"0de40008";
        when 11x"288" => o_wb_dat <= x"002f0c19";
        when 11x"289" => o_wb_dat <= x"c8200046";
        when 11x"28a" => o_wb_dat <= x"e9400000";
        when 11x"28b" => o_wb_dat <= x"01201410";
        when 11x"28c" => o_wb_dat <= x"01c01a10";
        when 11x"28d" => o_wb_dat <= x"00a01410";
        when 11x"28e" => o_wb_dat <= x"01001a10";
        when 11x"28f" => o_wb_dat <= x"00290c19";
        when 11x"290" => o_wb_dat <= x"c820001a";
        when 11x"291" => o_wb_dat <= x"c900003e";
        when 11x"292" => o_wb_dat <= x"89260003";
        when 11x"293" => o_wb_dat <= x"01400c10";
        when 11x"294" => o_wb_dat <= x"55c97ff8";
        when 11x"295" => o_wb_dat <= x"0028141b";
        when 11x"296" => o_wb_dat <= x"0ce40014";
        when 11x"297" => o_wb_dat <= x"c820002f";
        when 11x"298" => o_wb_dat <= x"54c60001";
        when 11x"299" => o_wb_dat <= x"2cc4000c";
        when 11x"29a" => o_wb_dat <= x"01071187";
        when 11x"29b" => o_wb_dat <= x"2ca80000";
        when 11x"29c" => o_wb_dat <= x"2d680004";
        when 11x"29d" => o_wb_dat <= x"c0a00032";
        when 11x"29e" => o_wb_dat <= x"02000a10";
        when 11x"29f" => o_wb_dat <= x"48420100";
        when 11x"2a0" => o_wb_dat <= x"c0400005";
        when 11x"2a1" => o_wb_dat <= x"e8400000";
        when 11x"2a2" => o_wb_dat <= x"00200a10";
        when 11x"2a3" => o_wb_dat <= x"f7c00000";
        when 11x"2a4" => o_wb_dat <= x"e7c00118";
        when 11x"2a5" => o_wb_dat <= x"00202010";
        when 11x"2a6" => o_wb_dat <= x"0e1c0004";
        when 11x"2a7" => o_wb_dat <= x"0fdc0000";
        when 11x"2a8" => o_wb_dat <= x"579c0008";
        when 11x"2a9" => o_wb_dat <= x"e3c00000";
        when 11x"2aa" => o_wb_dat <= x"c1200016";
        when 11x"2ab" => o_wb_dat <= x"54ea7ff8";
        when 11x"2ac" => o_wb_dat <= x"0c240014";
        when 11x"2ad" => o_wb_dat <= x"00e10e15";
        when 11x"2ae" => o_wb_dat <= x"0c270000";
        when 11x"2af" => o_wb_dat <= x"0ce70004";
        when 11x"2b0" => o_wb_dat <= x"00210e15";
        when 11x"2b1" => o_wb_dat <= x"00e6121b";
        when 11x"2b2" => o_wb_dat <= x"c8e00010";
        when 11x"2b3" => o_wb_dat <= x"0de40014";
        when 11x"2b4" => o_wb_dat <= x"00ef1403";
        when 11x"2b5" => o_wb_dat <= x"00e10e16";
        when 11x"2b6" => o_wb_dat <= x"01e7161c";
        when 11x"2b7" => o_wb_dat <= x"c9e00006";
        when 11x"2b8" => o_wb_dat <= x"01ee0e1a";
        when 11x"2b9" => o_wb_dat <= x"c9e00004";
        when 11x"2ba" => o_wb_dat <= x"01c00e10";
        when 11x"2bb" => o_wb_dat <= x"00a00210";
        when 11x"2bc" => o_wb_dat <= x"01001210";
        when 11x"2bd" => o_wb_dat <= x"55290001";
        when 11x"2be" => o_wb_dat <= x"554a0008";
        when 11x"2bf" => o_wb_dat <= x"e3ffffd0";
        when 11x"2c0" => o_wb_dat <= x"0c240000";
        when 11x"2c1" => o_wb_dat <= x"e3fffff0";
        when 11x"2c2" => o_wb_dat <= x"0ce40000";
        when 11x"2c3" => o_wb_dat <= x"0de40004";
        when 11x"2c4" => o_wb_dat <= x"00e71e15";
        when 11x"2c5" => o_wb_dat <= x"e3fffff0";
        when 11x"2c6" => o_wb_dat <= x"00271c03";
        when 11x"2c7" => o_wb_dat <= x"0027120b";
        when 11x"2c8" => o_wb_dat <= x"01271215";
        when 11x"2c9" => o_wb_dat <= x"00e71c15";
        when 11x"2ca" => o_wb_dat <= x"0ce70004";
        when 11x"2cb" => o_wb_dat <= x"2ce90004";
        when 11x"2cc" => o_wb_dat <= x"554a7fff";
        when 11x"2cd" => o_wb_dat <= x"01201c10";
        when 11x"2ce" => o_wb_dat <= x"e3ffffc6";
        when 11x"2cf" => o_wb_dat <= x"558c0001";
        when 11x"2d0" => o_wb_dat <= x"54840018";
        when 11x"2d1" => o_wb_dat <= x"e3ffffac";
        when 11x"2d2" => o_wb_dat <= x"00c00210";
        when 11x"2d3" => o_wb_dat <= x"0d1f75b4";
        when 11x"2d4" => o_wb_dat <= x"f4a7fffe";
        when 11x"2d5" => o_wb_dat <= x"54a505c0";
        when 11x"2d6" => o_wb_dat <= x"e8600000";
        when 11x"2d7" => o_wb_dat <= x"0028061b";
        when 11x"2d8" => o_wb_dat <= x"c8200020";
        when 11x"2d9" => o_wb_dat <= x"0c850000";
        when 11x"2da" => o_wb_dat <= x"e8400000";
        when 11x"2db" => o_wb_dat <= x"e3e00018";
        when 11x"2dc" => o_wb_dat <= x"0ce50008";
        when 11x"2dd" => o_wb_dat <= x"00270587";
        when 11x"2de" => o_wb_dat <= x"0ce10000";
        when 11x"2df" => o_wb_dat <= x"00e60e18";
        when 11x"2e0" => o_wb_dat <= x"c8e00012";
        when 11x"2e1" => o_wb_dat <= x"54847fff";
        when 11x"2e2" => o_wb_dat <= x"00a30615";
        when 11x"2e3" => o_wb_dat <= x"00650615";
        when 11x"2e4" => o_wb_dat <= x"f4a7fffe";
        when 11x"2e5" => o_wb_dat <= x"54a50574";
        when 11x"2e6" => o_wb_dat <= x"00650787";
        when 11x"2e7" => o_wb_dat <= x"2c83000c";
        when 11x"2e8" => o_wb_dat <= x"54210008";
        when 11x"2e9" => o_wb_dat <= x"0062081b";
        when 11x"2ea" => o_wb_dat <= x"c8600002";
        when 11x"2eb" => o_wb_dat <= x"e3c00000";
        when 11x"2ec" => o_wb_dat <= x"0c610000";
        when 11x"2ed" => o_wb_dat <= x"2c617ff8";
        when 11x"2ee" => o_wb_dat <= x"0ce10004";
        when 11x"2ef" => o_wb_dat <= x"2ce17ffc";
        when 11x"2f0" => o_wb_dat <= x"54420001";
        when 11x"2f1" => o_wb_dat <= x"e3fffff7";
        when 11x"2f2" => o_wb_dat <= x"54420001";
        when 11x"2f3" => o_wb_dat <= x"00220819";
        when 11x"2f4" => o_wb_dat <= x"c83fffe8";
        when 11x"2f5" => o_wb_dat <= x"54630001";
        when 11x"2f6" => o_wb_dat <= x"54a50018";
        when 11x"2f7" => o_wb_dat <= x"e3ffffe0";
        when 11x"2f8" => o_wb_dat <= x"e3c00000";
        when 11x"2f9" => o_wb_dat <= x"e820211c";
        when 11x"2fa" => o_wb_dat <= x"e3c00000";
        when 11x"2fb" => o_wb_dat <= x"579c7ffc";
        when 11x"2fc" => o_wb_dat <= x"2fdc0000";
        when 11x"2fd" => o_wb_dat <= x"ec580000";
        when 11x"2fe" => o_wb_dat <= x"0c620014";
        when 11x"2ff" => o_wb_dat <= x"0c820018";
        when 11x"300" => o_wb_dat <= x"ece80000";
        when 11x"301" => o_wb_dat <= x"2c270164";
        when 11x"302" => o_wb_dat <= x"54c1059c";
        when 11x"303" => o_wb_dat <= x"ece80000";
        when 11x"304" => o_wb_dat <= x"2cc7016c";
        when 11x"305" => o_wb_dat <= x"ece80000";
        when 11x"306" => o_wb_dat <= x"00c70c16";
        when 11x"307" => o_wb_dat <= x"8cc60002";
        when 11x"308" => o_wb_dat <= x"ed002800";
        when 11x"309" => o_wb_dat <= x"41080000";
        when 11x"30a" => o_wb_dat <= x"01080644";
        when 11x"30b" => o_wb_dat <= x"ecf04000";
        when 11x"30c" => o_wb_dat <= x"00e71010";
        when 11x"30d" => o_wb_dat <= x"2ce10000";
        when 11x"30e" => o_wb_dat <= x"ecf08000";
        when 11x"30f" => o_wb_dat <= x"00e70610";
        when 11x"310" => o_wb_dat <= x"2ce10004";
        when 11x"311" => o_wb_dat <= x"ecf0a000";
        when 11x"312" => o_wb_dat <= x"40e70005";
        when 11x"313" => o_wb_dat <= x"2ce10008";
        when 11x"314" => o_wb_dat <= x"ecec0000";
        when 11x"315" => o_wb_dat <= x"40e70001";
        when 11x"316" => o_wb_dat <= x"2ce1000c";
        when 11x"317" => o_wb_dat <= x"ecfff365";
        when 11x"318" => o_wb_dat <= x"40e7042e";
        when 11x"319" => o_wb_dat <= x"2ce10010";
        when 11x"31a" => o_wb_dat <= x"ecfffd6d";
        when 11x"31b" => o_wb_dat <= x"40e70570";
        when 11x"31c" => o_wb_dat <= x"2ce10014";
        when 11x"31d" => o_wb_dat <= x"54e10010";
        when 11x"31e" => o_wb_dat <= x"ed080000";
        when 11x"31f" => o_wb_dat <= x"2ce80168";
        when 11x"320" => o_wb_dat <= x"54210018";
        when 11x"321" => o_wb_dat <= x"ecf00000";
        when 11x"322" => o_wb_dat <= x"ed0a0000";
        when 11x"323" => o_wb_dat <= x"e96000b0";
        when 11x"324" => o_wb_dat <= x"e9200000";
        when 11x"325" => o_wb_dat <= x"01490841";
        when 11x"326" => o_wb_dat <= x"014a1644";
        when 11x"327" => o_wb_dat <= x"01481410";
        when 11x"328" => o_wb_dat <= x"2d410000";
        when 11x"329" => o_wb_dat <= x"55290001";
        when 11x"32a" => o_wb_dat <= x"01470c15";
        when 11x"32b" => o_wb_dat <= x"2d410004";
        when 11x"32c" => o_wb_dat <= x"54c6000a";
        when 11x"32d" => o_wb_dat <= x"54210008";
        when 11x"32e" => o_wb_dat <= x"5d4900b0";
        when 11x"32f" => o_wb_dat <= x"cd5ffff6";
        when 11x"330" => o_wb_dat <= x"ecea000f";
        when 11x"331" => o_wb_dat <= x"40e707ff";
        when 11x"332" => o_wb_dat <= x"2ce10000";
        when 11x"333" => o_wb_dat <= x"e7e0000c";
        when 11x"334" => o_wb_dat <= x"e7e00004";
        when 11x"335" => o_wb_dat <= x"0fdc0000";
        when 11x"336" => o_wb_dat <= x"579c0004";
        when 11x"337" => o_wb_dat <= x"e3c00000";
        when 11x"338" => o_wb_dat <= x"ec280000";
        when 11x"339" => o_wb_dat <= x"0c210164";
        when 11x"33a" => o_wb_dat <= x"ec480000";
        when 11x"33b" => o_wb_dat <= x"00220216";
        when 11x"33c" => o_wb_dat <= x"8c210002";
        when 11x"33d" => o_wb_dat <= x"2c220000";
        when 11x"33e" => o_wb_dat <= x"e3c00000";
        when 11x"33f" => o_wb_dat <= x"ec280000";
        when 11x"340" => o_wb_dat <= x"2c010170";
        when 11x"341" => o_wb_dat <= x"ec280000";
        when 11x"342" => o_wb_dat <= x"2c010174";
        when 11x"343" => o_wb_dat <= x"ec280000";
        when 11x"344" => o_wb_dat <= x"0c21016c";
        when 11x"345" => o_wb_dat <= x"e8400000";
        when 11x"346" => o_wb_dat <= x"e8601b80";
        when 11x"347" => o_wb_dat <= x"e3e00074";
        when 11x"348" => o_wb_dat <= x"ec680000";
        when 11x"349" => o_wb_dat <= x"0c630168";
        when 11x"34a" => o_wb_dat <= x"2c230000";
        when 11x"34b" => o_wb_dat <= x"2c430004";
        when 11x"34c" => o_wb_dat <= x"e3c00000";
        when 11x"34d" => o_wb_dat <= x"01403a10";
        when 11x"34e" => o_wb_dat <= x"ec400003";
        when 11x"34f" => o_wb_dat <= x"40420064";
        when 11x"350" => o_wb_dat <= x"ec680000";
        when 11x"351" => o_wb_dat <= x"0c630170";
        when 11x"352" => o_wb_dat <= x"ec880000";
        when 11x"353" => o_wb_dat <= x"0c840174";
        when 11x"354" => o_wb_dat <= x"ed080000";
        when 11x"355" => o_wb_dat <= x"0d08016c";
        when 11x"356" => o_wb_dat <= x"14a10000";
        when 11x"357" => o_wb_dat <= x"54210001";
        when 11x"358" => o_wb_dat <= x"c0a00033";
        when 11x"359" => o_wb_dat <= x"5cc5000a";
        when 11x"35a" => o_wb_dat <= x"c8c0001a";
        when 11x"35b" => o_wb_dat <= x"5cc5000d";
        when 11x"35c" => o_wb_dat <= x"ccc00003";
        when 11x"35d" => o_wb_dat <= x"e8600000";
        when 11x"35e" => o_wb_dat <= x"e3fffff8";
        when 11x"35f" => o_wb_dat <= x"5cc50009";
        when 11x"360" => o_wb_dat <= x"ccc00006";
        when 11x"361" => o_wb_dat <= x"54630008";
        when 11x"362" => o_wb_dat <= x"4c630007";
        when 11x"363" => o_wb_dat <= x"64c30028";
        when 11x"364" => o_wb_dat <= x"c8dffff2";
        when 11x"365" => o_wb_dat <= x"e3e0000f";
        when 11x"366" => o_wb_dat <= x"78a50020";
        when 11x"367" => o_wb_dat <= x"74a5007f";
        when 11x"368" => o_wb_dat <= x"54a57fe0";
        when 11x"369" => o_wb_dat <= x"00a20b87";
        when 11x"36a" => o_wb_dat <= x"eba00008";
        when 11x"36b" => o_wb_dat <= x"e8e00028";
        when 11x"36c" => o_wb_dat <= x"00c40e41";
        when 11x"36d" => o_wb_dat <= x"14258001";
        when 11x"36e" => o_wb_dat <= x"00c30d87";
        when 11x"36f" => o_wb_dat <= x"00c80c15";
        when 11x"370" => o_wb_dat <= x"00268e09";
        when 11x"371" => o_wb_dat <= x"54630001";
        when 11x"372" => o_wb_dat <= x"64a30028";
        when 11x"373" => o_wb_dat <= x"c8bfffe3";
        when 11x"374" => o_wb_dat <= x"e8600000";
        when 11x"375" => o_wb_dat <= x"54840001";
        when 11x"376" => o_wb_dat <= x"64a40016";
        when 11x"377" => o_wb_dat <= x"c8bfffdf";
        when 11x"378" => o_wb_dat <= x"e8800015";
        when 11x"379" => o_wb_dat <= x"54e80140";
        when 11x"37a" => o_wb_dat <= x"01201010";
        when 11x"37b" => o_wb_dat <= x"00a00000";
        when 11x"37c" => o_wb_dat <= x"e8c00690";
        when 11x"37d" => o_wb_dat <= x"03a50c1d";
        when 11x"37e" => o_wb_dat <= x"00dd0c16";
        when 11x"37f" => o_wb_dat <= x"0c278004";
        when 11x"380" => o_wb_dat <= x"00e73b07";
        when 11x"381" => o_wb_dat <= x"2c298004";
        when 11x"382" => o_wb_dat <= x"01293b07";
        when 11x"383" => o_wb_dat <= x"c4dffffa";
        when 11x"384" => o_wb_dat <= x"e8c00050";
        when 11x"385" => o_wb_dat <= x"03a50c1d";
        when 11x"386" => o_wb_dat <= x"00dd0c16";
        when 11x"387" => o_wb_dat <= x"2c098004";
        when 11x"388" => o_wb_dat <= x"01293b07";
        when 11x"389" => o_wb_dat <= x"c4dffffc";
        when 11x"38a" => o_wb_dat <= x"e3ffffcc";
        when 11x"38b" => o_wb_dat <= x"eca80000";
        when 11x"38c" => o_wb_dat <= x"2c650170";
        when 11x"38d" => o_wb_dat <= x"eca80000";
        when 11x"38e" => o_wb_dat <= x"2c850174";
        when 11x"38f" => o_wb_dat <= x"03a01410";
        when 11x"390" => o_wb_dat <= x"e3c00000";
        when 11x"391" => o_wb_dat <= x"579c7ff0";
        when 11x"392" => o_wb_dat <= x"2fdc000c";
        when 11x"393" => o_wb_dat <= x"ec800003";
        when 11x"394" => o_wb_dat <= x"40840052";
        when 11x"395" => o_wb_dat <= x"e8400008";
        when 11x"396" => o_wb_dat <= x"001c0409";
        when 11x"397" => o_wb_dat <= x"4861000f";
        when 11x"398" => o_wb_dat <= x"00640605";
        when 11x"399" => o_wb_dat <= x"54427fff";
        when 11x"39a" => o_wb_dat <= x"8c210004";
        when 11x"39b" => o_wb_dat <= x"007c0409";
        when 11x"39c" => o_wb_dat <= x"dc5ffffb";
        when 11x"39d" => o_wb_dat <= x"00203810";
        when 11x"39e" => o_wb_dat <= x"e7ffffaf";
        when 11x"39f" => o_wb_dat <= x"0fdc000c";
        when 11x"3a0" => o_wb_dat <= x"579c0010";
        when 11x"3a1" => o_wb_dat <= x"e3c00000";
        when 11x"3a2" => o_wb_dat <= x"579c7ff0";
        when 11x"3a3" => o_wb_dat <= x"2fdc000c";
        when 11x"3a4" => o_wb_dat <= x"ec800003";
        when 11x"3a5" => o_wb_dat <= x"40840052";
        when 11x"3a6" => o_wb_dat <= x"e840000b";
        when 11x"3a7" => o_wb_dat <= x"001c0409";
        when 11x"3a8" => o_wb_dat <= x"e8c0000a";
        when 11x"3a9" => o_wb_dat <= x"00a10019";
        when 11x"3aa" => o_wb_dat <= x"cca00002";
        when 11x"3ab" => o_wb_dat <= x"00210016";
        when 11x"3ac" => o_wb_dat <= x"00610c47";
        when 11x"3ad" => o_wb_dat <= x"54427fff";
        when 11x"3ae" => o_wb_dat <= x"00640605";
        when 11x"3af" => o_wb_dat <= x"00210c45";
        when 11x"3b0" => o_wb_dat <= x"007c0409";
        when 11x"3b1" => o_wb_dat <= x"c43ffffb";
        when 11x"3b2" => o_wb_dat <= x"cca00004";
        when 11x"3b3" => o_wb_dat <= x"e860002d";
        when 11x"3b4" => o_wb_dat <= x"54427fff";
        when 11x"3b5" => o_wb_dat <= x"007c0409";
        when 11x"3b6" => o_wb_dat <= x"003c0407";
        when 11x"3b7" => o_wb_dat <= x"e7ffff96";
        when 11x"3b8" => o_wb_dat <= x"0fdc000c";
        when 11x"3b9" => o_wb_dat <= x"579c0010";
        when 11x"3ba" => o_wb_dat <= x"e3c00000";
        when 11x"3bb" => o_wb_dat <= x"00c03a10";
        when 11x"3bc" => o_wb_dat <= x"c0600017";
        when 11x"3bd" => o_wb_dat <= x"00e00210";
        when 11x"3be" => o_wb_dat <= x"03a00000";
        when 11x"3bf" => o_wb_dat <= x"90420000";
        when 11x"3c0" => o_wb_dat <= x"00208410";
        when 11x"3c1" => o_wb_dat <= x"48a70003";
        when 11x"3c2" => o_wb_dat <= x"c0a00007";
        when 11x"3c3" => o_wb_dat <= x"58a50004";
        when 11x"3c4" => o_wb_dat <= x"03a30a1d";
        when 11x"3c5" => o_wb_dat <= x"007d0616";
        when 11x"3c6" => o_wb_dat <= x"24278001";
        when 11x"3c7" => o_wb_dat <= x"00e73a07";
        when 11x"3c8" => o_wb_dat <= x"c060000b";
        when 11x"3c9" => o_wb_dat <= x"00800000";
        when 11x"3ca" => o_wb_dat <= x"8ca30002";
        when 11x"3cb" => o_wb_dat <= x"c0a00006";
        when 11x"3cc" => o_wb_dat <= x"03a5081d";
        when 11x"3cd" => o_wb_dat <= x"00bd0a16";
        when 11x"3ce" => o_wb_dat <= x"2c278004";
        when 11x"3cf" => o_wb_dat <= x"00e73b07";
        when 11x"3d0" => o_wb_dat <= x"c4bffffc";
        when 11x"3d1" => o_wb_dat <= x"4ba30003";
        when 11x"3d2" => o_wb_dat <= x"24278001";
        when 11x"3d3" => o_wb_dat <= x"03a00c10";
        when 11x"3d4" => o_wb_dat <= x"e3c00000";
        when 11x"3d5" => o_wb_dat <= x"00c90000";
        when 11x"3d6" => o_wb_dat <= x"025b0192";
        when 11x"3d7" => o_wb_dat <= x"03ed0324";
        when 11x"3d8" => o_wb_dat <= x"057f04b6";
        when 11x"3d9" => o_wb_dat <= x"07110648";
        when 11x"3da" => o_wb_dat <= x"08a207d9";
        when 11x"3db" => o_wb_dat <= x"0a33096a";
        when 11x"3dc" => o_wb_dat <= x"0bc40afb";
        when 11x"3dd" => o_wb_dat <= x"0d540c8c";
        when 11x"3de" => o_wb_dat <= x"0ee30e1c";
        when 11x"3df" => o_wb_dat <= x"10720fab";
        when 11x"3e0" => o_wb_dat <= x"1201113a";
        when 11x"3e1" => o_wb_dat <= x"138f12c8";
        when 11x"3e2" => o_wb_dat <= x"151c1455";
        when 11x"3e3" => o_wb_dat <= x"16a815e2";
        when 11x"3e4" => o_wb_dat <= x"1833176e";
        when 11x"3e5" => o_wb_dat <= x"19be18f9";
        when 11x"3e6" => o_wb_dat <= x"1b471a82";
        when 11x"3e7" => o_wb_dat <= x"1ccf1c0b";
        when 11x"3e8" => o_wb_dat <= x"1e571d93";
        when 11x"3e9" => o_wb_dat <= x"1fdd1f1a";
        when 11x"3ea" => o_wb_dat <= x"2161209f";
        when 11x"3eb" => o_wb_dat <= x"22e52223";
        when 11x"3ec" => o_wb_dat <= x"246723a6";
        when 11x"3ed" => o_wb_dat <= x"25e82528";
        when 11x"3ee" => o_wb_dat <= x"276726a8";
        when 11x"3ef" => o_wb_dat <= x"28e52826";
        when 11x"3f0" => o_wb_dat <= x"2a6129a3";
        when 11x"3f1" => o_wb_dat <= x"2bdc2b1f";
        when 11x"3f2" => o_wb_dat <= x"2d552c99";
        when 11x"3f3" => o_wb_dat <= x"2ecc2e11";
        when 11x"3f4" => o_wb_dat <= x"30412f87";
        when 11x"3f5" => o_wb_dat <= x"31b530fb";
        when 11x"3f6" => o_wb_dat <= x"3326326e";
        when 11x"3f7" => o_wb_dat <= x"349633df";
        when 11x"3f8" => o_wb_dat <= x"3604354d";
        when 11x"3f9" => o_wb_dat <= x"376f36ba";
        when 11x"3fa" => o_wb_dat <= x"38d93824";
        when 11x"3fb" => o_wb_dat <= x"3a40398c";
        when 11x"3fc" => o_wb_dat <= x"3ba53af2";
        when 11x"3fd" => o_wb_dat <= x"3d073c56";
        when 11x"3fe" => o_wb_dat <= x"3e683db8";
        when 11x"3ff" => o_wb_dat <= x"3fc53f17";
        when 11x"400" => o_wb_dat <= x"41214073";
        when 11x"401" => o_wb_dat <= x"427a41ce";
        when 11x"402" => o_wb_dat <= x"43d04325";
        when 11x"403" => o_wb_dat <= x"4524447a";
        when 11x"404" => o_wb_dat <= x"467545cd";
        when 11x"405" => o_wb_dat <= x"47c3471c";
        when 11x"406" => o_wb_dat <= x"490f4869";
        when 11x"407" => o_wb_dat <= x"4a5849b4";
        when 11x"408" => o_wb_dat <= x"4b9d4afb";
        when 11x"409" => o_wb_dat <= x"4ce04c3f";
        when 11x"40a" => o_wb_dat <= x"4e204d81";
        when 11x"40b" => o_wb_dat <= x"4f5d4ebf";
        when 11x"40c" => o_wb_dat <= x"50974ffb";
        when 11x"40d" => o_wb_dat <= x"51ce5133";
        when 11x"40e" => o_wb_dat <= x"53025268";
        when 11x"40f" => o_wb_dat <= x"5432539b";
        when 11x"410" => o_wb_dat <= x"556054c9";
        when 11x"411" => o_wb_dat <= x"568a55f5";
        when 11x"412" => o_wb_dat <= x"57b0571d";
        when 11x"413" => o_wb_dat <= x"58d35842";
        when 11x"414" => o_wb_dat <= x"59f35964";
        when 11x"415" => o_wb_dat <= x"5b0f5a82";
        when 11x"416" => o_wb_dat <= x"5c285b9c";
        when 11x"417" => o_wb_dat <= x"5d3e5cb3";
        when 11x"418" => o_wb_dat <= x"5e4f5dc7";
        when 11x"419" => o_wb_dat <= x"5f5d5ed7";
        when 11x"41a" => o_wb_dat <= x"60685fe3";
        when 11x"41b" => o_wb_dat <= x"616e60eb";
        when 11x"41c" => o_wb_dat <= x"627161f0";
        when 11x"41d" => o_wb_dat <= x"637062f1";
        when 11x"41e" => o_wb_dat <= x"646c63ee";
        when 11x"41f" => o_wb_dat <= x"656364e8";
        when 11x"420" => o_wb_dat <= x"665665dd";
        when 11x"421" => o_wb_dat <= x"674666cf";
        when 11x"422" => o_wb_dat <= x"683267bc";
        when 11x"423" => o_wb_dat <= x"691968a6";
        when 11x"424" => o_wb_dat <= x"69fd698b";
        when 11x"425" => o_wb_dat <= x"6adc6a6d";
        when 11x"426" => o_wb_dat <= x"6bb76b4a";
        when 11x"427" => o_wb_dat <= x"6c8e6c23";
        when 11x"428" => o_wb_dat <= x"6d616cf8";
        when 11x"429" => o_wb_dat <= x"6e306dc9";
        when 11x"42a" => o_wb_dat <= x"6efb6e96";
        when 11x"42b" => o_wb_dat <= x"6fc16f5e";
        when 11x"42c" => o_wb_dat <= x"70837022";
        when 11x"42d" => o_wb_dat <= x"714070e2";
        when 11x"42e" => o_wb_dat <= x"71f9719d";
        when 11x"42f" => o_wb_dat <= x"72ae7254";
        when 11x"430" => o_wb_dat <= x"735e7307";
        when 11x"431" => o_wb_dat <= x"740a73b5";
        when 11x"432" => o_wb_dat <= x"74b2745f";
        when 11x"433" => o_wb_dat <= x"75557504";
        when 11x"434" => o_wb_dat <= x"75f375a5";
        when 11x"435" => o_wb_dat <= x"768d7641";
        when 11x"436" => o_wb_dat <= x"772276d8";
        when 11x"437" => o_wb_dat <= x"77b3776b";
        when 11x"438" => o_wb_dat <= x"783f77fa";
        when 11x"439" => o_wb_dat <= x"78c77884";
        when 11x"43a" => o_wb_dat <= x"794a7909";
        when 11x"43b" => o_wb_dat <= x"79c87989";
        when 11x"43c" => o_wb_dat <= x"7a417a05";
        when 11x"43d" => o_wb_dat <= x"7ab67a7c";
        when 11x"43e" => o_wb_dat <= x"7b267aee";
        when 11x"43f" => o_wb_dat <= x"7b917b5c";
        when 11x"440" => o_wb_dat <= x"7bf87bc5";
        when 11x"441" => o_wb_dat <= x"7c597c29";
        when 11x"442" => o_wb_dat <= x"7cb67c88";
        when 11x"443" => o_wb_dat <= x"7d0e7ce3";
        when 11x"444" => o_wb_dat <= x"7d627d39";
        when 11x"445" => o_wb_dat <= x"7db07d89";
        when 11x"446" => o_wb_dat <= x"7dfa7dd5";
        when 11x"447" => o_wb_dat <= x"7e3e7e1d";
        when 11x"448" => o_wb_dat <= x"7e7e7e5f";
        when 11x"449" => o_wb_dat <= x"7eb97e9c";
        when 11x"44a" => o_wb_dat <= x"7eef7ed5";
        when 11x"44b" => o_wb_dat <= x"7f217f09";
        when 11x"44c" => o_wb_dat <= x"7f4d7f37";
        when 11x"44d" => o_wb_dat <= x"7f747f61";
        when 11x"44e" => o_wb_dat <= x"7f977f86";
        when 11x"44f" => o_wb_dat <= x"7fb47fa6";
        when 11x"450" => o_wb_dat <= x"7fcd7fc1";
        when 11x"451" => o_wb_dat <= x"7fe17fd8";
        when 11x"452" => o_wb_dat <= x"7ff07fe9";
        when 11x"453" => o_wb_dat <= x"7ff97ff5";
        when 11x"454" => o_wb_dat <= x"7ffe7ffd";
        when 11x"455" => o_wb_dat <= x"7ffe7fff";
        when 11x"456" => o_wb_dat <= x"7ff97ffd";
        when 11x"457" => o_wb_dat <= x"7ff07ff5";
        when 11x"458" => o_wb_dat <= x"7fe17fe9";
        when 11x"459" => o_wb_dat <= x"7fcd7fd8";
        when 11x"45a" => o_wb_dat <= x"7fb47fc1";
        when 11x"45b" => o_wb_dat <= x"7f977fa6";
        when 11x"45c" => o_wb_dat <= x"7f747f86";
        when 11x"45d" => o_wb_dat <= x"7f4d7f61";
        when 11x"45e" => o_wb_dat <= x"7f217f37";
        when 11x"45f" => o_wb_dat <= x"7eef7f09";
        when 11x"460" => o_wb_dat <= x"7eb97ed5";
        when 11x"461" => o_wb_dat <= x"7e7e7e9c";
        when 11x"462" => o_wb_dat <= x"7e3e7e5f";
        when 11x"463" => o_wb_dat <= x"7dfa7e1d";
        when 11x"464" => o_wb_dat <= x"7db07dd5";
        when 11x"465" => o_wb_dat <= x"7d627d89";
        when 11x"466" => o_wb_dat <= x"7d0e7d39";
        when 11x"467" => o_wb_dat <= x"7cb67ce3";
        when 11x"468" => o_wb_dat <= x"7c597c88";
        when 11x"469" => o_wb_dat <= x"7bf87c29";
        when 11x"46a" => o_wb_dat <= x"7b917bc5";
        when 11x"46b" => o_wb_dat <= x"7b267b5c";
        when 11x"46c" => o_wb_dat <= x"7ab67aee";
        when 11x"46d" => o_wb_dat <= x"7a417a7c";
        when 11x"46e" => o_wb_dat <= x"79c87a05";
        when 11x"46f" => o_wb_dat <= x"794a7989";
        when 11x"470" => o_wb_dat <= x"78c77909";
        when 11x"471" => o_wb_dat <= x"783f7884";
        when 11x"472" => o_wb_dat <= x"77b377fa";
        when 11x"473" => o_wb_dat <= x"7722776b";
        when 11x"474" => o_wb_dat <= x"768d76d8";
        when 11x"475" => o_wb_dat <= x"75f37641";
        when 11x"476" => o_wb_dat <= x"755575a5";
        when 11x"477" => o_wb_dat <= x"74b27504";
        when 11x"478" => o_wb_dat <= x"740a745f";
        when 11x"479" => o_wb_dat <= x"735e73b5";
        when 11x"47a" => o_wb_dat <= x"72ae7307";
        when 11x"47b" => o_wb_dat <= x"71f97254";
        when 11x"47c" => o_wb_dat <= x"7140719d";
        when 11x"47d" => o_wb_dat <= x"708370e2";
        when 11x"47e" => o_wb_dat <= x"6fc17022";
        when 11x"47f" => o_wb_dat <= x"6efb6f5e";
        when 11x"480" => o_wb_dat <= x"6e306e96";
        when 11x"481" => o_wb_dat <= x"6d616dc9";
        when 11x"482" => o_wb_dat <= x"6c8e6cf8";
        when 11x"483" => o_wb_dat <= x"6bb76c23";
        when 11x"484" => o_wb_dat <= x"6adc6b4a";
        when 11x"485" => o_wb_dat <= x"69fd6a6d";
        when 11x"486" => o_wb_dat <= x"6919698b";
        when 11x"487" => o_wb_dat <= x"683268a6";
        when 11x"488" => o_wb_dat <= x"674667bc";
        when 11x"489" => o_wb_dat <= x"665666cf";
        when 11x"48a" => o_wb_dat <= x"656365dd";
        when 11x"48b" => o_wb_dat <= x"646c64e8";
        when 11x"48c" => o_wb_dat <= x"637063ee";
        when 11x"48d" => o_wb_dat <= x"627162f1";
        when 11x"48e" => o_wb_dat <= x"616e61f0";
        when 11x"48f" => o_wb_dat <= x"606860eb";
        when 11x"490" => o_wb_dat <= x"5f5d5fe3";
        when 11x"491" => o_wb_dat <= x"5e4f5ed7";
        when 11x"492" => o_wb_dat <= x"5d3e5dc7";
        when 11x"493" => o_wb_dat <= x"5c285cb3";
        when 11x"494" => o_wb_dat <= x"5b0f5b9c";
        when 11x"495" => o_wb_dat <= x"59f35a82";
        when 11x"496" => o_wb_dat <= x"58d35964";
        when 11x"497" => o_wb_dat <= x"57b05842";
        when 11x"498" => o_wb_dat <= x"568a571d";
        when 11x"499" => o_wb_dat <= x"556055f5";
        when 11x"49a" => o_wb_dat <= x"543254c9";
        when 11x"49b" => o_wb_dat <= x"5302539b";
        when 11x"49c" => o_wb_dat <= x"51ce5268";
        when 11x"49d" => o_wb_dat <= x"50975133";
        when 11x"49e" => o_wb_dat <= x"4f5d4ffb";
        when 11x"49f" => o_wb_dat <= x"4e204ebf";
        when 11x"4a0" => o_wb_dat <= x"4ce04d81";
        when 11x"4a1" => o_wb_dat <= x"4b9d4c3f";
        when 11x"4a2" => o_wb_dat <= x"4a584afb";
        when 11x"4a3" => o_wb_dat <= x"490f49b4";
        when 11x"4a4" => o_wb_dat <= x"47c34869";
        when 11x"4a5" => o_wb_dat <= x"4675471c";
        when 11x"4a6" => o_wb_dat <= x"452445cd";
        when 11x"4a7" => o_wb_dat <= x"43d0447a";
        when 11x"4a8" => o_wb_dat <= x"427a4325";
        when 11x"4a9" => o_wb_dat <= x"412141ce";
        when 11x"4aa" => o_wb_dat <= x"3fc54073";
        when 11x"4ab" => o_wb_dat <= x"3e683f17";
        when 11x"4ac" => o_wb_dat <= x"3d073db8";
        when 11x"4ad" => o_wb_dat <= x"3ba53c56";
        when 11x"4ae" => o_wb_dat <= x"3a403af2";
        when 11x"4af" => o_wb_dat <= x"38d9398c";
        when 11x"4b0" => o_wb_dat <= x"376f3824";
        when 11x"4b1" => o_wb_dat <= x"360436ba";
        when 11x"4b2" => o_wb_dat <= x"3496354d";
        when 11x"4b3" => o_wb_dat <= x"332633df";
        when 11x"4b4" => o_wb_dat <= x"31b5326e";
        when 11x"4b5" => o_wb_dat <= x"304130fb";
        when 11x"4b6" => o_wb_dat <= x"2ecc2f87";
        when 11x"4b7" => o_wb_dat <= x"2d552e11";
        when 11x"4b8" => o_wb_dat <= x"2bdc2c99";
        when 11x"4b9" => o_wb_dat <= x"2a612b1f";
        when 11x"4ba" => o_wb_dat <= x"28e529a3";
        when 11x"4bb" => o_wb_dat <= x"27672826";
        when 11x"4bc" => o_wb_dat <= x"25e826a8";
        when 11x"4bd" => o_wb_dat <= x"24672528";
        when 11x"4be" => o_wb_dat <= x"22e523a6";
        when 11x"4bf" => o_wb_dat <= x"21612223";
        when 11x"4c0" => o_wb_dat <= x"1fdd209f";
        when 11x"4c1" => o_wb_dat <= x"1e571f1a";
        when 11x"4c2" => o_wb_dat <= x"1ccf1d93";
        when 11x"4c3" => o_wb_dat <= x"1b471c0b";
        when 11x"4c4" => o_wb_dat <= x"19be1a82";
        when 11x"4c5" => o_wb_dat <= x"183318f9";
        when 11x"4c6" => o_wb_dat <= x"16a8176e";
        when 11x"4c7" => o_wb_dat <= x"151c15e2";
        when 11x"4c8" => o_wb_dat <= x"138f1455";
        when 11x"4c9" => o_wb_dat <= x"120112c8";
        when 11x"4ca" => o_wb_dat <= x"1072113a";
        when 11x"4cb" => o_wb_dat <= x"0ee30fab";
        when 11x"4cc" => o_wb_dat <= x"0d540e1c";
        when 11x"4cd" => o_wb_dat <= x"0bc40c8c";
        when 11x"4ce" => o_wb_dat <= x"0a330afb";
        when 11x"4cf" => o_wb_dat <= x"08a2096a";
        when 11x"4d0" => o_wb_dat <= x"071107d9";
        when 11x"4d1" => o_wb_dat <= x"057f0648";
        when 11x"4d2" => o_wb_dat <= x"03ed04b6";
        when 11x"4d3" => o_wb_dat <= x"025b0324";
        when 11x"4d4" => o_wb_dat <= x"00c90192";
        when 11x"4d5" => o_wb_dat <= x"ff370000";
        when 11x"4d6" => o_wb_dat <= x"fda5fe6e";
        when 11x"4d7" => o_wb_dat <= x"fc13fcdc";
        when 11x"4d8" => o_wb_dat <= x"fa81fb4a";
        when 11x"4d9" => o_wb_dat <= x"f8eff9b8";
        when 11x"4da" => o_wb_dat <= x"f75ef827";
        when 11x"4db" => o_wb_dat <= x"f5cdf696";
        when 11x"4dc" => o_wb_dat <= x"f43cf505";
        when 11x"4dd" => o_wb_dat <= x"f2acf374";
        when 11x"4de" => o_wb_dat <= x"f11df1e4";
        when 11x"4df" => o_wb_dat <= x"ef8ef055";
        when 11x"4e0" => o_wb_dat <= x"edffeec6";
        when 11x"4e1" => o_wb_dat <= x"ec71ed38";
        when 11x"4e2" => o_wb_dat <= x"eae4ebab";
        when 11x"4e3" => o_wb_dat <= x"e958ea1e";
        when 11x"4e4" => o_wb_dat <= x"e7cde892";
        when 11x"4e5" => o_wb_dat <= x"e642e707";
        when 11x"4e6" => o_wb_dat <= x"e4b9e57e";
        when 11x"4e7" => o_wb_dat <= x"e331e3f5";
        when 11x"4e8" => o_wb_dat <= x"e1a9e26d";
        when 11x"4e9" => o_wb_dat <= x"e023e0e6";
        when 11x"4ea" => o_wb_dat <= x"de9fdf61";
        when 11x"4eb" => o_wb_dat <= x"dd1bdddd";
        when 11x"4ec" => o_wb_dat <= x"db99dc5a";
        when 11x"4ed" => o_wb_dat <= x"da18dad8";
        when 11x"4ee" => o_wb_dat <= x"d899d958";
        when 11x"4ef" => o_wb_dat <= x"d71bd7da";
        when 11x"4f0" => o_wb_dat <= x"d59fd65d";
        when 11x"4f1" => o_wb_dat <= x"d424d4e1";
        when 11x"4f2" => o_wb_dat <= x"d2abd367";
        when 11x"4f3" => o_wb_dat <= x"d134d1ef";
        when 11x"4f4" => o_wb_dat <= x"cfbfd079";
        when 11x"4f5" => o_wb_dat <= x"ce4bcf05";
        when 11x"4f6" => o_wb_dat <= x"ccdacd92";
        when 11x"4f7" => o_wb_dat <= x"cb6acc21";
        when 11x"4f8" => o_wb_dat <= x"c9fccab3";
        when 11x"4f9" => o_wb_dat <= x"c891c946";
        when 11x"4fa" => o_wb_dat <= x"c727c7dc";
        when 11x"4fb" => o_wb_dat <= x"c5c0c674";
        when 11x"4fc" => o_wb_dat <= x"c45bc50e";
        when 11x"4fd" => o_wb_dat <= x"c2f9c3aa";
        when 11x"4fe" => o_wb_dat <= x"c198c248";
        when 11x"4ff" => o_wb_dat <= x"c03bc0e9";
        when 11x"500" => o_wb_dat <= x"bedfbf8d";
        when 11x"501" => o_wb_dat <= x"bd86be32";
        when 11x"502" => o_wb_dat <= x"bc30bcdb";
        when 11x"503" => o_wb_dat <= x"badcbb86";
        when 11x"504" => o_wb_dat <= x"b98bba33";
        when 11x"505" => o_wb_dat <= x"b83db8e4";
        when 11x"506" => o_wb_dat <= x"b6f1b797";
        when 11x"507" => o_wb_dat <= x"b5a8b64c";
        when 11x"508" => o_wb_dat <= x"b463b505";
        when 11x"509" => o_wb_dat <= x"b320b3c1";
        when 11x"50a" => o_wb_dat <= x"b1e0b27f";
        when 11x"50b" => o_wb_dat <= x"b0a3b141";
        when 11x"50c" => o_wb_dat <= x"af69b005";
        when 11x"50d" => o_wb_dat <= x"ae32aecd";
        when 11x"50e" => o_wb_dat <= x"acfead98";
        when 11x"50f" => o_wb_dat <= x"abceac65";
        when 11x"510" => o_wb_dat <= x"aaa0ab37";
        when 11x"511" => o_wb_dat <= x"a976aa0b";
        when 11x"512" => o_wb_dat <= x"a850a8e3";
        when 11x"513" => o_wb_dat <= x"a72da7be";
        when 11x"514" => o_wb_dat <= x"a60da69c";
        when 11x"515" => o_wb_dat <= x"a4f1a57e";
        when 11x"516" => o_wb_dat <= x"a3d8a464";
        when 11x"517" => o_wb_dat <= x"a2c2a34d";
        when 11x"518" => o_wb_dat <= x"a1b1a239";
        when 11x"519" => o_wb_dat <= x"a0a3a129";
        when 11x"51a" => o_wb_dat <= x"9f98a01d";
        when 11x"51b" => o_wb_dat <= x"9e929f15";
        when 11x"51c" => o_wb_dat <= x"9d8f9e10";
        when 11x"51d" => o_wb_dat <= x"9c909d0f";
        when 11x"51e" => o_wb_dat <= x"9b949c12";
        when 11x"51f" => o_wb_dat <= x"9a9d9b18";
        when 11x"520" => o_wb_dat <= x"99aa9a23";
        when 11x"521" => o_wb_dat <= x"98ba9931";
        when 11x"522" => o_wb_dat <= x"97ce9844";
        when 11x"523" => o_wb_dat <= x"96e7975a";
        when 11x"524" => o_wb_dat <= x"96039675";
        when 11x"525" => o_wb_dat <= x"95249593";
        when 11x"526" => o_wb_dat <= x"944994b6";
        when 11x"527" => o_wb_dat <= x"937293dd";
        when 11x"528" => o_wb_dat <= x"929f9308";
        when 11x"529" => o_wb_dat <= x"91d09237";
        when 11x"52a" => o_wb_dat <= x"9105916a";
        when 11x"52b" => o_wb_dat <= x"903f90a2";
        when 11x"52c" => o_wb_dat <= x"8f7d8fde";
        when 11x"52d" => o_wb_dat <= x"8ec08f1e";
        when 11x"52e" => o_wb_dat <= x"8e078e63";
        when 11x"52f" => o_wb_dat <= x"8d528dac";
        when 11x"530" => o_wb_dat <= x"8ca28cf9";
        when 11x"531" => o_wb_dat <= x"8bf68c4b";
        when 11x"532" => o_wb_dat <= x"8b4e8ba1";
        when 11x"533" => o_wb_dat <= x"8aab8afc";
        when 11x"534" => o_wb_dat <= x"8a0d8a5b";
        when 11x"535" => o_wb_dat <= x"897389bf";
        when 11x"536" => o_wb_dat <= x"88de8928";
        when 11x"537" => o_wb_dat <= x"884d8895";
        when 11x"538" => o_wb_dat <= x"87c18806";
        when 11x"539" => o_wb_dat <= x"8739877c";
        when 11x"53a" => o_wb_dat <= x"86b686f7";
        when 11x"53b" => o_wb_dat <= x"86388677";
        when 11x"53c" => o_wb_dat <= x"85bf85fb";
        when 11x"53d" => o_wb_dat <= x"854a8584";
        when 11x"53e" => o_wb_dat <= x"84da8512";
        when 11x"53f" => o_wb_dat <= x"846f84a4";
        when 11x"540" => o_wb_dat <= x"8408843b";
        when 11x"541" => o_wb_dat <= x"83a783d7";
        when 11x"542" => o_wb_dat <= x"834a8378";
        when 11x"543" => o_wb_dat <= x"82f2831d";
        when 11x"544" => o_wb_dat <= x"829e82c7";
        when 11x"545" => o_wb_dat <= x"82508277";
        when 11x"546" => o_wb_dat <= x"8206822b";
        when 11x"547" => o_wb_dat <= x"81c281e3";
        when 11x"548" => o_wb_dat <= x"818281a1";
        when 11x"549" => o_wb_dat <= x"81478164";
        when 11x"54a" => o_wb_dat <= x"8111812b";
        when 11x"54b" => o_wb_dat <= x"80df80f7";
        when 11x"54c" => o_wb_dat <= x"80b380c9";
        when 11x"54d" => o_wb_dat <= x"808c809f";
        when 11x"54e" => o_wb_dat <= x"8069807a";
        when 11x"54f" => o_wb_dat <= x"804c805a";
        when 11x"550" => o_wb_dat <= x"8033803f";
        when 11x"551" => o_wb_dat <= x"801f8028";
        when 11x"552" => o_wb_dat <= x"80108017";
        when 11x"553" => o_wb_dat <= x"8007800b";
        when 11x"554" => o_wb_dat <= x"80028003";
        when 11x"555" => o_wb_dat <= x"80028001";
        when 11x"556" => o_wb_dat <= x"80078003";
        when 11x"557" => o_wb_dat <= x"8010800b";
        when 11x"558" => o_wb_dat <= x"801f8017";
        when 11x"559" => o_wb_dat <= x"80338028";
        when 11x"55a" => o_wb_dat <= x"804c803f";
        when 11x"55b" => o_wb_dat <= x"8069805a";
        when 11x"55c" => o_wb_dat <= x"808c807a";
        when 11x"55d" => o_wb_dat <= x"80b3809f";
        when 11x"55e" => o_wb_dat <= x"80df80c9";
        when 11x"55f" => o_wb_dat <= x"811180f7";
        when 11x"560" => o_wb_dat <= x"8147812b";
        when 11x"561" => o_wb_dat <= x"81828164";
        when 11x"562" => o_wb_dat <= x"81c281a1";
        when 11x"563" => o_wb_dat <= x"820681e3";
        when 11x"564" => o_wb_dat <= x"8250822b";
        when 11x"565" => o_wb_dat <= x"829e8277";
        when 11x"566" => o_wb_dat <= x"82f282c7";
        when 11x"567" => o_wb_dat <= x"834a831d";
        when 11x"568" => o_wb_dat <= x"83a78378";
        when 11x"569" => o_wb_dat <= x"840883d7";
        when 11x"56a" => o_wb_dat <= x"846f843b";
        when 11x"56b" => o_wb_dat <= x"84da84a4";
        when 11x"56c" => o_wb_dat <= x"854a8512";
        when 11x"56d" => o_wb_dat <= x"85bf8584";
        when 11x"56e" => o_wb_dat <= x"863885fb";
        when 11x"56f" => o_wb_dat <= x"86b68677";
        when 11x"570" => o_wb_dat <= x"873986f7";
        when 11x"571" => o_wb_dat <= x"87c1877c";
        when 11x"572" => o_wb_dat <= x"884d8806";
        when 11x"573" => o_wb_dat <= x"88de8895";
        when 11x"574" => o_wb_dat <= x"89738928";
        when 11x"575" => o_wb_dat <= x"8a0d89bf";
        when 11x"576" => o_wb_dat <= x"8aab8a5b";
        when 11x"577" => o_wb_dat <= x"8b4e8afc";
        when 11x"578" => o_wb_dat <= x"8bf68ba1";
        when 11x"579" => o_wb_dat <= x"8ca28c4b";
        when 11x"57a" => o_wb_dat <= x"8d528cf9";
        when 11x"57b" => o_wb_dat <= x"8e078dac";
        when 11x"57c" => o_wb_dat <= x"8ec08e63";
        when 11x"57d" => o_wb_dat <= x"8f7d8f1e";
        when 11x"57e" => o_wb_dat <= x"903f8fde";
        when 11x"57f" => o_wb_dat <= x"910590a2";
        when 11x"580" => o_wb_dat <= x"91d0916a";
        when 11x"581" => o_wb_dat <= x"929f9237";
        when 11x"582" => o_wb_dat <= x"93729308";
        when 11x"583" => o_wb_dat <= x"944993dd";
        when 11x"584" => o_wb_dat <= x"952494b6";
        when 11x"585" => o_wb_dat <= x"96039593";
        when 11x"586" => o_wb_dat <= x"96e79675";
        when 11x"587" => o_wb_dat <= x"97ce975a";
        when 11x"588" => o_wb_dat <= x"98ba9844";
        when 11x"589" => o_wb_dat <= x"99aa9931";
        when 11x"58a" => o_wb_dat <= x"9a9d9a23";
        when 11x"58b" => o_wb_dat <= x"9b949b18";
        when 11x"58c" => o_wb_dat <= x"9c909c12";
        when 11x"58d" => o_wb_dat <= x"9d8f9d0f";
        when 11x"58e" => o_wb_dat <= x"9e929e10";
        when 11x"58f" => o_wb_dat <= x"9f989f15";
        when 11x"590" => o_wb_dat <= x"a0a3a01d";
        when 11x"591" => o_wb_dat <= x"a1b1a129";
        when 11x"592" => o_wb_dat <= x"a2c2a239";
        when 11x"593" => o_wb_dat <= x"a3d8a34d";
        when 11x"594" => o_wb_dat <= x"a4f1a464";
        when 11x"595" => o_wb_dat <= x"a60da57e";
        when 11x"596" => o_wb_dat <= x"a72da69c";
        when 11x"597" => o_wb_dat <= x"a850a7be";
        when 11x"598" => o_wb_dat <= x"a976a8e3";
        when 11x"599" => o_wb_dat <= x"aaa0aa0b";
        when 11x"59a" => o_wb_dat <= x"abceab37";
        when 11x"59b" => o_wb_dat <= x"acfeac65";
        when 11x"59c" => o_wb_dat <= x"ae32ad98";
        when 11x"59d" => o_wb_dat <= x"af69aecd";
        when 11x"59e" => o_wb_dat <= x"b0a3b005";
        when 11x"59f" => o_wb_dat <= x"b1e0b141";
        when 11x"5a0" => o_wb_dat <= x"b320b27f";
        when 11x"5a1" => o_wb_dat <= x"b463b3c1";
        when 11x"5a2" => o_wb_dat <= x"b5a8b505";
        when 11x"5a3" => o_wb_dat <= x"b6f1b64c";
        when 11x"5a4" => o_wb_dat <= x"b83db797";
        when 11x"5a5" => o_wb_dat <= x"b98bb8e4";
        when 11x"5a6" => o_wb_dat <= x"badcba33";
        when 11x"5a7" => o_wb_dat <= x"bc30bb86";
        when 11x"5a8" => o_wb_dat <= x"bd86bcdb";
        when 11x"5a9" => o_wb_dat <= x"bedfbe32";
        when 11x"5aa" => o_wb_dat <= x"c03bbf8d";
        when 11x"5ab" => o_wb_dat <= x"c198c0e9";
        when 11x"5ac" => o_wb_dat <= x"c2f9c248";
        when 11x"5ad" => o_wb_dat <= x"c45bc3aa";
        when 11x"5ae" => o_wb_dat <= x"c5c0c50e";
        when 11x"5af" => o_wb_dat <= x"c727c674";
        when 11x"5b0" => o_wb_dat <= x"c891c7dc";
        when 11x"5b1" => o_wb_dat <= x"c9fcc946";
        when 11x"5b2" => o_wb_dat <= x"cb6acab3";
        when 11x"5b3" => o_wb_dat <= x"ccdacc21";
        when 11x"5b4" => o_wb_dat <= x"ce4bcd92";
        when 11x"5b5" => o_wb_dat <= x"cfbfcf05";
        when 11x"5b6" => o_wb_dat <= x"d134d079";
        when 11x"5b7" => o_wb_dat <= x"d2abd1ef";
        when 11x"5b8" => o_wb_dat <= x"d424d367";
        when 11x"5b9" => o_wb_dat <= x"d59fd4e1";
        when 11x"5ba" => o_wb_dat <= x"d71bd65d";
        when 11x"5bb" => o_wb_dat <= x"d899d7da";
        when 11x"5bc" => o_wb_dat <= x"da18d958";
        when 11x"5bd" => o_wb_dat <= x"db99dad8";
        when 11x"5be" => o_wb_dat <= x"dd1bdc5a";
        when 11x"5bf" => o_wb_dat <= x"de9fdddd";
        when 11x"5c0" => o_wb_dat <= x"e023df61";
        when 11x"5c1" => o_wb_dat <= x"e1a9e0e6";
        when 11x"5c2" => o_wb_dat <= x"e331e26d";
        when 11x"5c3" => o_wb_dat <= x"e4b9e3f5";
        when 11x"5c4" => o_wb_dat <= x"e642e57e";
        when 11x"5c5" => o_wb_dat <= x"e7cde707";
        when 11x"5c6" => o_wb_dat <= x"e958e892";
        when 11x"5c7" => o_wb_dat <= x"eae4ea1e";
        when 11x"5c8" => o_wb_dat <= x"ec71ebab";
        when 11x"5c9" => o_wb_dat <= x"edffed38";
        when 11x"5ca" => o_wb_dat <= x"ef8eeec6";
        when 11x"5cb" => o_wb_dat <= x"f11df055";
        when 11x"5cc" => o_wb_dat <= x"f2acf1e4";
        when 11x"5cd" => o_wb_dat <= x"f43cf374";
        when 11x"5ce" => o_wb_dat <= x"f5cdf505";
        when 11x"5cf" => o_wb_dat <= x"f75ef696";
        when 11x"5d0" => o_wb_dat <= x"f8eff827";
        when 11x"5d1" => o_wb_dat <= x"fa81f9b8";
        when 11x"5d2" => o_wb_dat <= x"fc13fb4a";
        when 11x"5d3" => o_wb_dat <= x"fda5fcdc";
        when 11x"5d4" => o_wb_dat <= x"ff37fe6e";
        when 11x"5d5" => o_wb_dat <= x"00001758";
        when 11x"5d6" => o_wb_dat <= x"676f7270";
        when 11x"5d7" => o_wb_dat <= x"006d6172";
        when 11x"5d8" => o_wb_dat <= x"2031434d";
        when 11x"5d9" => o_wb_dat <= x"6854202d";
        when 11x"5da" => o_wb_dat <= x"524d2065";
        when 11x"5db" => o_wb_dat <= x"33435349";
        when 11x"5dc" => o_wb_dat <= x"6f632032";
        when 11x"5dd" => o_wb_dat <= x"7475706d";
        when 11x"5de" => o_wb_dat <= x"0a0a7265";
        when 11x"5df" => o_wb_dat <= x"41525600";
        when 11x"5e0" => o_wb_dat <= x"20203a4d";
        when 11x"5e1" => o_wb_dat <= x"58007830";
        when 11x"5e2" => o_wb_dat <= x"3a4d4152";
        when 11x"5e3" => o_wb_dat <= x"78302020";
        when 11x"5e4" => o_wb_dat <= x"53534200";
        when 11x"5e5" => o_wb_dat <= x"2020203a";
        when 11x"5e6" => o_wb_dat <= x"56007830";
        when 11x"5e7" => o_wb_dat <= x"3a4e4f43";
        when 11x"5e8" => o_wb_dat <= x"78302020";
        when 11x"5e9" => o_wb_dat <= x"61745300";
        when 11x"5ea" => o_wb_dat <= x"203a6b63";
        when 11x"5eb" => o_wb_dat <= x"2c007830";
        when 11x"5ec" => o_wb_dat <= x"62200020";
        when 11x"5ed" => o_wb_dat <= x"73657479";
        when 11x"5ee" => o_wb_dat <= x"410a000a";
        when 11x"5ef" => o_wb_dat <= x"45444342";
        when 11x"5f0" => o_wb_dat <= x"49484746";
        when 11x"5f1" => o_wb_dat <= x"4d4c4b4a";
        when 11x"5f2" => o_wb_dat <= x"51504f4e";
        when 11x"5f3" => o_wb_dat <= x"55545352";
        when 11x"5f4" => o_wb_dat <= x"59585756";
        when 11x"5f5" => o_wb_dat <= x"62610a5a";
        when 11x"5f6" => o_wb_dat <= x"66656463";
        when 11x"5f7" => o_wb_dat <= x"6a696867";
        when 11x"5f8" => o_wb_dat <= x"6e6d6c6b";
        when 11x"5f9" => o_wb_dat <= x"7271706f";
        when 11x"5fa" => o_wb_dat <= x"76757473";
        when 11x"5fb" => o_wb_dat <= x"7a797877";
        when 11x"5fc" => o_wb_dat <= x"3231300a";
        when 11x"5fd" => o_wb_dat <= x"36353433";
        when 11x"5fe" => o_wb_dat <= x"0a393837";
        when 11x"5ff" => o_wb_dat <= x"3f212e2c";
        when 11x"600" => o_wb_dat <= x"25242322";
        when 11x"601" => o_wb_dat <= x"5b292826";
        when 11x"602" => o_wb_dat <= x"3c7d7b5d";
        when 11x"603" => o_wb_dat <= x"2d2b3d3e";
        when 11x"604" => o_wb_dat <= x"5c7c2f2a";
        when 11x"605" => o_wb_dat <= x"09410a7e";
        when 11x"606" => o_wb_dat <= x"09430942";
        when 11x"607" => o_wb_dat <= x"00000a44";
        when 11x"608" => o_wb_dat <= x"6f6d654d";
        when 11x"609" => o_wb_dat <= x"70207972";
        when 11x"60a" => o_wb_dat <= x"3a6c6f6f";
        when 11x"60b" => o_wb_dat <= x"3020200a";
        when 11x"60c" => o_wb_dat <= x"00000078";
        when 11x"60d" => o_wb_dat <= x"0000202c";
        when 11x"60e" => o_wb_dat <= x"74796220";
        when 11x"60f" => o_wb_dat <= x"66207365";
        when 11x"610" => o_wb_dat <= x"0a656572";
        when 11x"611" => o_wb_dat <= x"79542020";
        when 11x"612" => o_wb_dat <= x"203a6570";
        when 11x"613" => o_wb_dat <= x"00000000";
        when 11x"614" => o_wb_dat <= x"3130000a";
        when 11x"615" => o_wb_dat <= x"35343332";
        when 11x"616" => o_wb_dat <= x"39383736";
        when 11x"617" => o_wb_dat <= x"44434241";
        when 11x"618" => o_wb_dat <= x"00004645";
        when 11x"619" => o_wb_dat <= x"00000000";
        when 11x"61a" => o_wb_dat <= x"00000000";
        when 11x"61b" => o_wb_dat <= x"08080808";
        when 11x"61c" => o_wb_dat <= x"00080008";
        when 11x"61d" => o_wb_dat <= x"00001414";
        when 11x"61e" => o_wb_dat <= x"00000000";
        when 11x"61f" => o_wb_dat <= x"22227f22";
        when 11x"620" => o_wb_dat <= x"00227f22";
        when 11x"621" => o_wb_dat <= x"3e017e14";
        when 11x"622" => o_wb_dat <= x"00143f40";
        when 11x"623" => o_wb_dat <= x"08122542";
        when 11x"624" => o_wb_dat <= x"00215224";
        when 11x"625" => o_wb_dat <= x"040a120c";
        when 11x"626" => o_wb_dat <= x"006e112a";
        when 11x"627" => o_wb_dat <= x"00000808";
        when 11x"628" => o_wb_dat <= x"00000000";
        when 11x"629" => o_wb_dat <= x"04040810";
        when 11x"62a" => o_wb_dat <= x"00100804";
        when 11x"62b" => o_wb_dat <= x"10100804";
        when 11x"62c" => o_wb_dat <= x"00040810";
        when 11x"62d" => o_wb_dat <= x"1c2a0800";
        when 11x"62e" => o_wb_dat <= x"00002214";
        when 11x"62f" => o_wb_dat <= x"3e080800";
        when 11x"630" => o_wb_dat <= x"00000808";
        when 11x"631" => o_wb_dat <= x"00000000";
        when 11x"632" => o_wb_dat <= x"00040800";
        when 11x"633" => o_wb_dat <= x"3e000000";
        when 11x"634" => o_wb_dat <= x"00000000";
        when 11x"635" => o_wb_dat <= x"00000000";
        when 11x"636" => o_wb_dat <= x"00080000";
        when 11x"637" => o_wb_dat <= x"08102040";
        when 11x"638" => o_wb_dat <= x"00010204";
        when 11x"639" => o_wb_dat <= x"4951613e";
        when 11x"63a" => o_wb_dat <= x"003e4345";
        when 11x"63b" => o_wb_dat <= x"08080c08";
        when 11x"63c" => o_wb_dat <= x"001c0808";
        when 11x"63d" => o_wb_dat <= x"1820413e";
        when 11x"63e" => o_wb_dat <= x"007f0204";
        when 11x"63f" => o_wb_dat <= x"3c40413e";
        when 11x"640" => o_wb_dat <= x"003e4140";
        when 11x"641" => o_wb_dat <= x"22242830";
        when 11x"642" => o_wb_dat <= x"0020207f";
        when 11x"643" => o_wb_dat <= x"3f01017f";
        when 11x"644" => o_wb_dat <= x"003e4140";
        when 11x"645" => o_wb_dat <= x"3f01021c";
        when 11x"646" => o_wb_dat <= x"003e4141";
        when 11x"647" => o_wb_dat <= x"1020407f";
        when 11x"648" => o_wb_dat <= x"00040408";
        when 11x"649" => o_wb_dat <= x"3e41413e";
        when 11x"64a" => o_wb_dat <= x"003e4141";
        when 11x"64b" => o_wb_dat <= x"7e41413e";
        when 11x"64c" => o_wb_dat <= x"001c2040";
        when 11x"64d" => o_wb_dat <= x"00080000";
        when 11x"64e" => o_wb_dat <= x"00000800";
        when 11x"64f" => o_wb_dat <= x"00080000";
        when 11x"650" => o_wb_dat <= x"00040800";
        when 11x"651" => o_wb_dat <= x"02040810";
        when 11x"652" => o_wb_dat <= x"00100804";
        when 11x"653" => o_wb_dat <= x"007f0000";
        when 11x"654" => o_wb_dat <= x"0000007f";
        when 11x"655" => o_wb_dat <= x"20100804";
        when 11x"656" => o_wb_dat <= x"00040810";
        when 11x"657" => o_wb_dat <= x"3040413e";
        when 11x"658" => o_wb_dat <= x"00080008";
        when 11x"659" => o_wb_dat <= x"255d413e";
        when 11x"65a" => o_wb_dat <= x"003e411d";
        when 11x"65b" => o_wb_dat <= x"22221408";
        when 11x"65c" => o_wb_dat <= x"0041413e";
        when 11x"65d" => o_wb_dat <= x"3f41413f";
        when 11x"65e" => o_wb_dat <= x"003f4141";
        when 11x"65f" => o_wb_dat <= x"0101413e";
        when 11x"660" => o_wb_dat <= x"003e4101";
        when 11x"661" => o_wb_dat <= x"4141211f";
        when 11x"662" => o_wb_dat <= x"001f2141";
        when 11x"663" => o_wb_dat <= x"0f01017f";
        when 11x"664" => o_wb_dat <= x"007f0101";
        when 11x"665" => o_wb_dat <= x"0f01017f";
        when 11x"666" => o_wb_dat <= x"00010101";
        when 11x"667" => o_wb_dat <= x"7901413e";
        when 11x"668" => o_wb_dat <= x"003e4141";
        when 11x"669" => o_wb_dat <= x"7f414141";
        when 11x"66a" => o_wb_dat <= x"00414141";
        when 11x"66b" => o_wb_dat <= x"0808081c";
        when 11x"66c" => o_wb_dat <= x"001c0808";
        when 11x"66d" => o_wb_dat <= x"20202020";
        when 11x"66e" => o_wb_dat <= x"001c2220";
        when 11x"66f" => o_wb_dat <= x"0f112141";
        when 11x"670" => o_wb_dat <= x"00412111";
        when 11x"671" => o_wb_dat <= x"01010101";
        when 11x"672" => o_wb_dat <= x"007f0101";
        when 11x"673" => o_wb_dat <= x"49556341";
        when 11x"674" => o_wb_dat <= x"00414141";
        when 11x"675" => o_wb_dat <= x"49454341";
        when 11x"676" => o_wb_dat <= x"00416151";
        when 11x"677" => o_wb_dat <= x"4141221c";
        when 11x"678" => o_wb_dat <= x"001c2241";
        when 11x"679" => o_wb_dat <= x"3f41413f";
        when 11x"67a" => o_wb_dat <= x"00010101";
        when 11x"67b" => o_wb_dat <= x"4141221c";
        when 11x"67c" => o_wb_dat <= x"005c2251";
        when 11x"67d" => o_wb_dat <= x"3f41413f";
        when 11x"67e" => o_wb_dat <= x"00412111";
        when 11x"67f" => o_wb_dat <= x"3e01413e";
        when 11x"680" => o_wb_dat <= x"003e4140";
        when 11x"681" => o_wb_dat <= x"0808087f";
        when 11x"682" => o_wb_dat <= x"00080808";
        when 11x"683" => o_wb_dat <= x"41414141";
        when 11x"684" => o_wb_dat <= x"003e4141";
        when 11x"685" => o_wb_dat <= x"22414141";
        when 11x"686" => o_wb_dat <= x"00081422";
        when 11x"687" => o_wb_dat <= x"49414141";
        when 11x"688" => o_wb_dat <= x"00416355";
        when 11x"689" => o_wb_dat <= x"08142241";
        when 11x"68a" => o_wb_dat <= x"00412214";
        when 11x"68b" => o_wb_dat <= x"08142241";
        when 11x"68c" => o_wb_dat <= x"00080808";
        when 11x"68d" => o_wb_dat <= x"3e10207f";
        when 11x"68e" => o_wb_dat <= x"007f0204";
        when 11x"68f" => o_wb_dat <= x"0404041c";
        when 11x"690" => o_wb_dat <= x"001c0404";
        when 11x"691" => o_wb_dat <= x"08040201";
        when 11x"692" => o_wb_dat <= x"00402010";
        when 11x"693" => o_wb_dat <= x"1010101c";
        when 11x"694" => o_wb_dat <= x"001c1010";
        when 11x"695" => o_wb_dat <= x"00001408";
        when 11x"696" => o_wb_dat <= x"00000000";
        when 11x"697" => o_wb_dat <= x"00000000";
        when 11x"698" => o_wb_dat <= x"007f0000";
        when 11x"699" => o_wb_dat <= x"00000804";
        when 11x"69a" => o_wb_dat <= x"00000000";
        when 11x"69b" => o_wb_dat <= x"201e0000";
        when 11x"69c" => o_wb_dat <= x"005e213e";
        when 11x"69d" => o_wb_dat <= x"463a0202";
        when 11x"69e" => o_wb_dat <= x"003d4242";
        when 11x"69f" => o_wb_dat <= x"013e0000";
        when 11x"6a0" => o_wb_dat <= x"003e0101";
        when 11x"6a1" => o_wb_dat <= x"312e2020";
        when 11x"6a2" => o_wb_dat <= x"005e2121";
        when 11x"6a3" => o_wb_dat <= x"211e0000";
        when 11x"6a4" => o_wb_dat <= x"001e013f";
        when 11x"6a5" => o_wb_dat <= x"0e041408";
        when 11x"6a6" => o_wb_dat <= x"00040404";
        when 11x"6a7" => o_wb_dat <= x"213e0000";
        when 11x"6a8" => o_wb_dat <= x"1e203e21";
        when 11x"6a9" => o_wb_dat <= x"231d0101";
        when 11x"6aa" => o_wb_dat <= x"00212121";
        when 11x"6ab" => o_wb_dat <= x"08000800";
        when 11x"6ac" => o_wb_dat <= x"00080808";
        when 11x"6ad" => o_wb_dat <= x"08000800";
        when 11x"6ae" => o_wb_dat <= x"06080808";
        when 11x"6af" => o_wb_dat <= x"09110101";
        when 11x"6b0" => o_wb_dat <= x"00110907";
        when 11x"6b1" => o_wb_dat <= x"04040404";
        when 11x"6b2" => o_wb_dat <= x"00080404";
        when 11x"6b3" => o_wb_dat <= x"4b350000";
        when 11x"6b4" => o_wb_dat <= x"00494949";
        when 11x"6b5" => o_wb_dat <= x"231d0000";
        when 11x"6b6" => o_wb_dat <= x"00212121";
        when 11x"6b7" => o_wb_dat <= x"211e0000";
        when 11x"6b8" => o_wb_dat <= x"001e2121";
        when 11x"6b9" => o_wb_dat <= x"221e0000";
        when 11x"6ba" => o_wb_dat <= x"02021e22";
        when 11x"6bb" => o_wb_dat <= x"223c0000";
        when 11x"6bc" => o_wb_dat <= x"20203c22";
        when 11x"6bd" => o_wb_dat <= x"231d0000";
        when 11x"6be" => o_wb_dat <= x"00010101";
        when 11x"6bf" => o_wb_dat <= x"023c0000";
        when 11x"6c0" => o_wb_dat <= x"001e201c";
        when 11x"6c1" => o_wb_dat <= x"040e0400";
        when 11x"6c2" => o_wb_dat <= x"00180404";
        when 11x"6c3" => o_wb_dat <= x"22220000";
        when 11x"6c4" => o_wb_dat <= x"005c2222";
        when 11x"6c5" => o_wb_dat <= x"22220000";
        when 11x"6c6" => o_wb_dat <= x"00081414";
        when 11x"6c7" => o_wb_dat <= x"41410000";
        when 11x"6c8" => o_wb_dat <= x"00225549";
        when 11x"6c9" => o_wb_dat <= x"14220000";
        when 11x"6ca" => o_wb_dat <= x"00221408";
        when 11x"6cb" => o_wb_dat <= x"22220000";
        when 11x"6cc" => o_wb_dat <= x"1c202c32";
        when 11x"6cd" => o_wb_dat <= x"203e0000";
        when 11x"6ce" => o_wb_dat <= x"003e0408";
        when 11x"6cf" => o_wb_dat <= x"02040418";
        when 11x"6d0" => o_wb_dat <= x"00180404";
        when 11x"6d1" => o_wb_dat <= x"08080808";
        when 11x"6d2" => o_wb_dat <= x"00080808";
        when 11x"6d3" => o_wb_dat <= x"2010100c";
        when 11x"6d4" => o_wb_dat <= x"000c1010";
        when 11x"6d5" => o_wb_dat <= x"4c000000";
        when 11x"6d6" => o_wb_dat <= x"00000032";
        when 11x"6d7" => o_wb_dat <= x"00220000";
        when 11x"6d8" => o_wb_dat <= x"001c2200";
        when 11x"6d9" => o_wb_dat <= x"00000000";
        when 11x"6da" => o_wb_dat <= x"00000000";
        when 11x"6db" => o_wb_dat <= x"00000000";
        when 11x"6dc" => o_wb_dat <= x"00000000";
        when 11x"6dd" => o_wb_dat <= x"00000000";
        when 11x"6de" => o_wb_dat <= x"00000000";
        when 11x"6df" => o_wb_dat <= x"00000000";
        when 11x"6e0" => o_wb_dat <= x"00000000";
        when 11x"6e1" => o_wb_dat <= x"00000000";
        when 11x"6e2" => o_wb_dat <= x"00000000";
        when 11x"6e3" => o_wb_dat <= x"00000000";
        when 11x"6e4" => o_wb_dat <= x"00000000";
        when 11x"6e5" => o_wb_dat <= x"00000000";
        when 11x"6e6" => o_wb_dat <= x"00000000";
        when 11x"6e7" => o_wb_dat <= x"00000000";
        when 11x"6e8" => o_wb_dat <= x"00000000";
        when 11x"6e9" => o_wb_dat <= x"00000000";
        when 11x"6ea" => o_wb_dat <= x"00000000";
        when 11x"6eb" => o_wb_dat <= x"00000000";
        when 11x"6ec" => o_wb_dat <= x"00000000";
        when 11x"6ed" => o_wb_dat <= x"00000000";
        when 11x"6ee" => o_wb_dat <= x"00000000";
        when 11x"6ef" => o_wb_dat <= x"00000000";
        when 11x"6f0" => o_wb_dat <= x"00000000";
        when 11x"6f1" => o_wb_dat <= x"00000000";
        when 11x"6f2" => o_wb_dat <= x"00000000";
        when 11x"6f3" => o_wb_dat <= x"00000000";
        when 11x"6f4" => o_wb_dat <= x"00000000";
        when 11x"6f5" => o_wb_dat <= x"00000000";
        when 11x"6f6" => o_wb_dat <= x"00000000";
        when 11x"6f7" => o_wb_dat <= x"00000000";
        when 11x"6f8" => o_wb_dat <= x"00000000";
        when 11x"6f9" => o_wb_dat <= x"00000000";
        when 11x"6fa" => o_wb_dat <= x"00000000";
        when 11x"6fb" => o_wb_dat <= x"00000000";
        when 11x"6fc" => o_wb_dat <= x"00000000";
        when 11x"6fd" => o_wb_dat <= x"00000000";
        when 11x"6fe" => o_wb_dat <= x"00000000";
        when 11x"6ff" => o_wb_dat <= x"00000000";
        when 11x"700" => o_wb_dat <= x"00000000";
        when 11x"701" => o_wb_dat <= x"00000000";
        when 11x"702" => o_wb_dat <= x"00000000";
        when 11x"703" => o_wb_dat <= x"00000000";
        when 11x"704" => o_wb_dat <= x"00000000";
        when 11x"705" => o_wb_dat <= x"00000000";
        when 11x"706" => o_wb_dat <= x"00000000";
        when 11x"707" => o_wb_dat <= x"00000000";
        when 11x"708" => o_wb_dat <= x"00000000";
        when 11x"709" => o_wb_dat <= x"00000000";
        when 11x"70a" => o_wb_dat <= x"00000000";
        when 11x"70b" => o_wb_dat <= x"00000000";
        when 11x"70c" => o_wb_dat <= x"00000000";
        when 11x"70d" => o_wb_dat <= x"00000000";
        when 11x"70e" => o_wb_dat <= x"00000000";
        when 11x"70f" => o_wb_dat <= x"00000000";
        when 11x"710" => o_wb_dat <= x"00000000";
        when 11x"711" => o_wb_dat <= x"00000000";
        when 11x"712" => o_wb_dat <= x"00000000";
        when 11x"713" => o_wb_dat <= x"00000000";
        when 11x"714" => o_wb_dat <= x"00000000";
        when 11x"715" => o_wb_dat <= x"00000000";
        when 11x"716" => o_wb_dat <= x"00000000";
        when 11x"717" => o_wb_dat <= x"00000000";
        when 11x"718" => o_wb_dat <= x"00000000";
        when 11x"719" => o_wb_dat <= x"00000000";
        when 11x"71a" => o_wb_dat <= x"00000000";
        when 11x"71b" => o_wb_dat <= x"00000000";
        when 11x"71c" => o_wb_dat <= x"00000000";
        when 11x"71d" => o_wb_dat <= x"00000000";
        when 11x"71e" => o_wb_dat <= x"00000000";
        when 11x"71f" => o_wb_dat <= x"00000000";
        when 11x"720" => o_wb_dat <= x"00000000";
        when 11x"721" => o_wb_dat <= x"00000000";
        when 11x"722" => o_wb_dat <= x"00000000";
        when 11x"723" => o_wb_dat <= x"00000000";
        when 11x"724" => o_wb_dat <= x"00000000";
        when 11x"725" => o_wb_dat <= x"00000000";
        when 11x"726" => o_wb_dat <= x"00000000";
        when 11x"727" => o_wb_dat <= x"00000000";
        when 11x"728" => o_wb_dat <= x"00000000";
        when 11x"729" => o_wb_dat <= x"00000000";
        when 11x"72a" => o_wb_dat <= x"00000000";
        when 11x"72b" => o_wb_dat <= x"00000000";
        when 11x"72c" => o_wb_dat <= x"00000000";
        when 11x"72d" => o_wb_dat <= x"00000000";
        when 11x"72e" => o_wb_dat <= x"00000000";
        when 11x"72f" => o_wb_dat <= x"00000000";
        when 11x"730" => o_wb_dat <= x"00000000";
        when 11x"731" => o_wb_dat <= x"00000000";
        when 11x"732" => o_wb_dat <= x"00000000";
        when 11x"733" => o_wb_dat <= x"00000000";
        when 11x"734" => o_wb_dat <= x"00000000";
        when 11x"735" => o_wb_dat <= x"00000000";
        when 11x"736" => o_wb_dat <= x"00000000";
        when 11x"737" => o_wb_dat <= x"00000000";
        when 11x"738" => o_wb_dat <= x"00000000";
        when 11x"739" => o_wb_dat <= x"00000000";
        when 11x"73a" => o_wb_dat <= x"00000000";
        when 11x"73b" => o_wb_dat <= x"00000000";
        when 11x"73c" => o_wb_dat <= x"00000000";
        when 11x"73d" => o_wb_dat <= x"00000000";
        when 11x"73e" => o_wb_dat <= x"00000000";
        when 11x"73f" => o_wb_dat <= x"00000000";
        when 11x"740" => o_wb_dat <= x"00000000";
        when 11x"741" => o_wb_dat <= x"00000000";
        when 11x"742" => o_wb_dat <= x"00000000";
        when 11x"743" => o_wb_dat <= x"00000000";
        when 11x"744" => o_wb_dat <= x"00000000";
        when 11x"745" => o_wb_dat <= x"00000000";
        when 11x"746" => o_wb_dat <= x"00000000";
        when 11x"747" => o_wb_dat <= x"00000000";
        when 11x"748" => o_wb_dat <= x"00000000";
        when 11x"749" => o_wb_dat <= x"00000000";
        when 11x"74a" => o_wb_dat <= x"00000000";
        when 11x"74b" => o_wb_dat <= x"00000000";
        when 11x"74c" => o_wb_dat <= x"00000000";
        when 11x"74d" => o_wb_dat <= x"00000000";
        when 11x"74e" => o_wb_dat <= x"00000000";
        when 11x"74f" => o_wb_dat <= x"00000000";
        when 11x"750" => o_wb_dat <= x"00000000";
        when 11x"751" => o_wb_dat <= x"00000000";
        when 11x"752" => o_wb_dat <= x"00000000";
        when 11x"753" => o_wb_dat <= x"00000000";
        when 11x"754" => o_wb_dat <= x"00000000";
        when 11x"755" => o_wb_dat <= x"00000000";
        when 11x"756" => o_wb_dat <= x"00000000";
        when 11x"757" => o_wb_dat <= x"00000000";
        when 11x"758" => o_wb_dat <= x"00000000";
        when 11x"759" => o_wb_dat <= x"00000000";
        when 11x"75a" => o_wb_dat <= x"00000000";
        when 11x"75b" => o_wb_dat <= x"00000000";
        when 11x"75c" => o_wb_dat <= x"00000000";
        when 11x"75d" => o_wb_dat <= x"00000000";
        when 11x"75e" => o_wb_dat <= x"00000000";
        when 11x"75f" => o_wb_dat <= x"00000000";
        when 11x"760" => o_wb_dat <= x"00000000";
        when 11x"761" => o_wb_dat <= x"00000000";
        when 11x"762" => o_wb_dat <= x"00000000";
        when 11x"763" => o_wb_dat <= x"00000000";
        when 11x"764" => o_wb_dat <= x"00000000";
        when 11x"765" => o_wb_dat <= x"00000000";
        when 11x"766" => o_wb_dat <= x"00000000";
        when 11x"767" => o_wb_dat <= x"00000000";
        when 11x"768" => o_wb_dat <= x"00000000";
        when 11x"769" => o_wb_dat <= x"00000000";
        when 11x"76a" => o_wb_dat <= x"00000000";
        when 11x"76b" => o_wb_dat <= x"00000000";
        when 11x"76c" => o_wb_dat <= x"00000000";
        when 11x"76d" => o_wb_dat <= x"00000000";
        when 11x"76e" => o_wb_dat <= x"00000000";
        when 11x"76f" => o_wb_dat <= x"00000000";
        when 11x"770" => o_wb_dat <= x"00000000";
        when 11x"771" => o_wb_dat <= x"00000000";
        when 11x"772" => o_wb_dat <= x"00000000";
        when 11x"773" => o_wb_dat <= x"00000000";
        when 11x"774" => o_wb_dat <= x"00000000";
        when 11x"775" => o_wb_dat <= x"00000000";
        when 11x"776" => o_wb_dat <= x"00000000";
        when 11x"777" => o_wb_dat <= x"00000000";
        when 11x"778" => o_wb_dat <= x"00000000";
        when 11x"779" => o_wb_dat <= x"00000000";
        when 11x"77a" => o_wb_dat <= x"00000000";
        when 11x"77b" => o_wb_dat <= x"00000000";
        when 11x"77c" => o_wb_dat <= x"00000000";
        when 11x"77d" => o_wb_dat <= x"00000000";
        when 11x"77e" => o_wb_dat <= x"00000000";
        when 11x"77f" => o_wb_dat <= x"00000000";
        when 11x"780" => o_wb_dat <= x"00000000";
        when 11x"781" => o_wb_dat <= x"00000000";
        when 11x"782" => o_wb_dat <= x"00000000";
        when 11x"783" => o_wb_dat <= x"00000000";
        when 11x"784" => o_wb_dat <= x"00000000";
        when 11x"785" => o_wb_dat <= x"00000000";
        when 11x"786" => o_wb_dat <= x"00000000";
        when 11x"787" => o_wb_dat <= x"00000000";
        when 11x"788" => o_wb_dat <= x"00000000";
        when 11x"789" => o_wb_dat <= x"00000000";
        when 11x"78a" => o_wb_dat <= x"00000000";
        when 11x"78b" => o_wb_dat <= x"00000000";
        when 11x"78c" => o_wb_dat <= x"00000000";
        when 11x"78d" => o_wb_dat <= x"00000000";
        when 11x"78e" => o_wb_dat <= x"00000000";
        when 11x"78f" => o_wb_dat <= x"00000000";
        when 11x"790" => o_wb_dat <= x"00000000";
        when 11x"791" => o_wb_dat <= x"00000000";
        when 11x"792" => o_wb_dat <= x"00000000";
        when 11x"793" => o_wb_dat <= x"00000000";
        when 11x"794" => o_wb_dat <= x"00000000";
        when 11x"795" => o_wb_dat <= x"00000000";
        when 11x"796" => o_wb_dat <= x"00000000";
        when 11x"797" => o_wb_dat <= x"00000000";
        when 11x"798" => o_wb_dat <= x"00000000";
        when 11x"799" => o_wb_dat <= x"00000000";
        when 11x"79a" => o_wb_dat <= x"00000000";
        when 11x"79b" => o_wb_dat <= x"00000000";
        when 11x"79c" => o_wb_dat <= x"00000000";
        when 11x"79d" => o_wb_dat <= x"00000000";
        when 11x"79e" => o_wb_dat <= x"00000000";
        when 11x"79f" => o_wb_dat <= x"00000000";
        when 11x"7a0" => o_wb_dat <= x"00000000";
        when 11x"7a1" => o_wb_dat <= x"00000000";
        when 11x"7a2" => o_wb_dat <= x"00000000";
        when 11x"7a3" => o_wb_dat <= x"00000000";
        when 11x"7a4" => o_wb_dat <= x"00000000";
        when 11x"7a5" => o_wb_dat <= x"00000000";
        when 11x"7a6" => o_wb_dat <= x"00000000";
        when 11x"7a7" => o_wb_dat <= x"00000000";
        when 11x"7a8" => o_wb_dat <= x"00000000";
        when 11x"7a9" => o_wb_dat <= x"00000000";
        when 11x"7aa" => o_wb_dat <= x"00000000";
        when 11x"7ab" => o_wb_dat <= x"00000000";
        when 11x"7ac" => o_wb_dat <= x"00000000";
        when 11x"7ad" => o_wb_dat <= x"00000000";
        when 11x"7ae" => o_wb_dat <= x"00000000";
        when 11x"7af" => o_wb_dat <= x"00000000";
        when 11x"7b0" => o_wb_dat <= x"00000000";
        when 11x"7b1" => o_wb_dat <= x"00000000";
        when 11x"7b2" => o_wb_dat <= x"00000000";
        when 11x"7b3" => o_wb_dat <= x"00000000";
        when 11x"7b4" => o_wb_dat <= x"00000000";
        when 11x"7b5" => o_wb_dat <= x"00000000";
        when 11x"7b6" => o_wb_dat <= x"00000000";
        when 11x"7b7" => o_wb_dat <= x"00000000";
        when 11x"7b8" => o_wb_dat <= x"00000000";
        when 11x"7b9" => o_wb_dat <= x"00000000";
        when 11x"7ba" => o_wb_dat <= x"00000000";
        when 11x"7bb" => o_wb_dat <= x"00000000";
        when 11x"7bc" => o_wb_dat <= x"00000000";
        when 11x"7bd" => o_wb_dat <= x"00000000";
        when 11x"7be" => o_wb_dat <= x"00000000";
        when 11x"7bf" => o_wb_dat <= x"00000000";
        when 11x"7c0" => o_wb_dat <= x"00000000";
        when 11x"7c1" => o_wb_dat <= x"00000000";
        when 11x"7c2" => o_wb_dat <= x"00000000";
        when 11x"7c3" => o_wb_dat <= x"00000000";
        when 11x"7c4" => o_wb_dat <= x"00000000";
        when 11x"7c5" => o_wb_dat <= x"00000000";
        when 11x"7c6" => o_wb_dat <= x"00000000";
        when 11x"7c7" => o_wb_dat <= x"00000000";
        when 11x"7c8" => o_wb_dat <= x"00000000";
        when 11x"7c9" => o_wb_dat <= x"00000000";
        when 11x"7ca" => o_wb_dat <= x"00000000";
        when 11x"7cb" => o_wb_dat <= x"00000000";
        when 11x"7cc" => o_wb_dat <= x"00000000";
        when 11x"7cd" => o_wb_dat <= x"00000000";
        when 11x"7ce" => o_wb_dat <= x"00000000";
        when 11x"7cf" => o_wb_dat <= x"00000000";
        when 11x"7d0" => o_wb_dat <= x"00000000";
        when 11x"7d1" => o_wb_dat <= x"00000000";
        when 11x"7d2" => o_wb_dat <= x"00000000";
        when 11x"7d3" => o_wb_dat <= x"00000000";
        when 11x"7d4" => o_wb_dat <= x"00000000";
        when 11x"7d5" => o_wb_dat <= x"00000000";
        when 11x"7d6" => o_wb_dat <= x"00000000";
        when 11x"7d7" => o_wb_dat <= x"00000000";
        when 11x"7d8" => o_wb_dat <= x"00000000";
        when 11x"7d9" => o_wb_dat <= x"00000000";
        when 11x"7da" => o_wb_dat <= x"00000000";
        when 11x"7db" => o_wb_dat <= x"00000000";
        when 11x"7dc" => o_wb_dat <= x"00000000";
        when 11x"7dd" => o_wb_dat <= x"00000000";
        when 11x"7de" => o_wb_dat <= x"00000000";
        when 11x"7df" => o_wb_dat <= x"00000000";
        when 11x"7e0" => o_wb_dat <= x"00000000";
        when 11x"7e1" => o_wb_dat <= x"00000000";
        when 11x"7e2" => o_wb_dat <= x"00000000";
        when 11x"7e3" => o_wb_dat <= x"00000000";
        when 11x"7e4" => o_wb_dat <= x"00000000";
        when 11x"7e5" => o_wb_dat <= x"00000000";
        when 11x"7e6" => o_wb_dat <= x"00000000";
        when 11x"7e7" => o_wb_dat <= x"00000000";
        when 11x"7e8" => o_wb_dat <= x"00000000";
        when 11x"7e9" => o_wb_dat <= x"00000000";
        when 11x"7ea" => o_wb_dat <= x"00000000";
        when 11x"7eb" => o_wb_dat <= x"00000000";
        when 11x"7ec" => o_wb_dat <= x"00000000";
        when 11x"7ed" => o_wb_dat <= x"00000000";
        when 11x"7ee" => o_wb_dat <= x"00000000";
        when 11x"7ef" => o_wb_dat <= x"00000000";
        when 11x"7f0" => o_wb_dat <= x"00000000";
        when 11x"7f1" => o_wb_dat <= x"00000000";
        when 11x"7f2" => o_wb_dat <= x"00000000";
        when 11x"7f3" => o_wb_dat <= x"00000000";
        when 11x"7f4" => o_wb_dat <= x"00000000";
        when 11x"7f5" => o_wb_dat <= x"00000000";
        when 11x"7f6" => o_wb_dat <= x"00000000";
        when 11x"7f7" => o_wb_dat <= x"00000000";
        when 11x"7f8" => o_wb_dat <= x"00000000";
        when 11x"7f9" => o_wb_dat <= x"00000000";
        when 11x"7fa" => o_wb_dat <= x"00000000";
        when 11x"7fb" => o_wb_dat <= x"00000000";
        when 11x"7fc" => o_wb_dat <= x"00000000";
        when 11x"7fd" => o_wb_dat <= x"00000000";
        when 11x"7fe" => o_wb_dat <= x"00000000";
        when 11x"7ff" => o_wb_dat <= x"00000000";

        when others => o_wb_dat <= (others => '0');
      end case;
    end if;
  end process;
end rtl;
