----------------------------------------------------------------------------------------------------
-- Copyright (c) 2019 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- This file contains common types for the video logic.
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package vid_types is
  --------------------------------------------------------------------------------------------------
  -- Video control registers.
  --------------------------------------------------------------------------------------------------
  type T_VID_REGS is record
    ADDR : std_logic_vector(23 downto 0);
    XOFFS : std_logic_vector(23 downto 0);
    XINCR : std_logic_vector(23 downto 0);
    HSTRT : std_logic_vector(23 downto 0);
    HSTOP : std_logic_vector(23 downto 0);
    CMODE : std_logic_vector(23 downto 0);
  end record T_VID_REGS;
end package;
