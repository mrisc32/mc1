----------------------------------------------------------------------------------------------------
-- Copyright (c) 2019 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- This is a single-ported ROM (Wishbone B4 pipelined interface).
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
  port(
    -- Control signals.
    i_clk : in std_logic;

    -- Wishbone memory interface (b4 pipelined slave).
    -- See: https://cdn.opencores.org/downloads/wbspec_b4.pdf
    i_wb_cyc : in std_logic;
    i_wb_stb : in std_logic;
    i_wb_adr : in std_logic_vector(31 downto 2);
    o_wb_dat : out std_logic_vector(31 downto 0);
    o_wb_ack : out std_logic;
    o_wb_stall : out std_logic
  );
end rom;

architecture rtl of rom is
  constant C_ADDR_BITS : positive := 9;
  constant C_ROM_SIZE : positive := 2**C_ADDR_BITS;

  type T_ROM_ARRAY is array (0 to C_ROM_SIZE-1) of std_logic_vector(31 downto 0);
  constant C_ROM_ARRAY : T_ROM_ARRAY := (
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"e8200000",
    x"e8400000",
    x"e8600000",
    x"e8800000",
    x"e8a00000",
    x"e8c00000",
    x"e8e00000",
    x"e9000000",
    x"e9200000",
    x"e9400000",
    x"e9600000",
    x"e9800000",
    x"e9a00000",
    x"e9c00000",
    x"e9e00000",
    x"ea000000",
    x"ea200000",
    x"ea400000",
    x"ea600000",
    x"ea800000",
    x"eaa00000",
    x"eac00000",
    x"eae00000",
    x"eb000000",
    x"eb200000",
    x"eb400000",
    x"eb600000",
    x"eb800000",
    x"eba00000",
    x"ebc00000",
    x"03a00000",
    x"40208000",
    x"40408000",
    x"40608000",
    x"40808000",
    x"40a08000",
    x"40c08000",
    x"40e08000",
    x"41008000",
    x"41208000",
    x"41408000",
    x"41608000",
    x"41808000",
    x"41a08000",
    x"41c08000",
    x"41e08000",
    x"42008000",
    x"42208000",
    x"42408000",
    x"42608000",
    x"42808000",
    x"42a08000",
    x"42c08000",
    x"42e08000",
    x"43008000",
    x"43208000",
    x"43408000",
    x"43608000",
    x"43808000",
    x"43a08000",
    x"43c08000",
    x"43e08000",
    x"eba00000",
    x"40208000",
    x"40408000",
    x"40608000",
    x"40808000",
    x"40a08000",
    x"40c08000",
    x"40e08000",
    x"41008000",
    x"41208000",
    x"41408000",
    x"41608000",
    x"41808000",
    x"41a08000",
    x"41c08000",
    x"41e08000",
    x"42008000",
    x"42208000",
    x"42408000",
    x"42608000",
    x"42808000",
    x"42a08000",
    x"42c08000",
    x"42e08000",
    x"43008000",
    x"43208000",
    x"43408000",
    x"43608000",
    x"43808000",
    x"43a08000",
    x"43c08000",
    x"43e08000",
    x"03a00000",
    x"ef880080",
    x"579c0000",
    x"e8200001",
    x"ec400000",
    x"544206b4",
    x"ede00000",
    x"e5e000f1",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"e3e00000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"579c7ffc",
    x"2fdc0000",
    x"e7e00005",
    x"e7e00064",
    x"0fdc0000",
    x"579c0004",
    x"e3c00000",
    x"579c7ffc",
    x"2fbc0000",
    x"ed680000",
    x"416b0000",
    x"ed904010",
    x"2d8b0000",
    x"ed90a000",
    x"418c0002",
    x"2d8b0004",
    x"ed90c000",
    x"418c0001",
    x"2d8b0008",
    x"ed8c0000",
    x"418c00ff",
    x"2d8b000c",
    x"556b0010",
    x"e8200064",
    x"e8400032",
    x"e8600000",
    x"e8800002",
    x"e8a00003",
    x"e8c00001",
    x"edffe000",
    x"2deb0000",
    x"e9c00001",
    x"88e30010",
    x"89020008",
    x"00e71010",
    x"00e70210",
    x"00e71e10",
    x"00eb1d0b",
    x"00210815",
    x"6ce100ff",
    x"0100021b",
    x"00e71012",
    x"c8e00003",
    x"00840016",
    x"00210815",
    x"00420a15",
    x"6ce200ff",
    x"0100041b",
    x"00e71012",
    x"c8e00003",
    x"00a50016",
    x"00420a15",
    x"00630c15",
    x"6ce300ff",
    x"0100061b",
    x"00e71012",
    x"c8e00003",
    x"00c60016",
    x"00630c15",
    x"55ce0001",
    x"60ee0100",
    x"c8ffffe3",
    x"556b0400",
    x"ec2a0000",
    x"ec500000",
    x"40420400",
    x"2c2b0000",
    x"2c4b0004",
    x"ed908000",
    x"418c0500",
    x"2d8b0008",
    x"556b000c",
    x"e3e00004",
    x"2c2b0000",
    x"2c4b0004",
    x"556b0008",
    x"54210002",
    x"544200a0",
    x"49a13fff",
    x"65ad02d0",
    x"c9bffff9",
    x"ed8a000f",
    x"418c07ff",
    x"2d8b0000",
    x"ed280002",
    x"41290000",
    x"01400000",
    x"e960e100",
    x"03aa161d",
    x"017d1616",
    x"2c098004",
    x"01293b07",
    x"c57ffffc",
    x"0fbc0000",
    x"579c0004",
    x"e3c00000",
    x"d8200006",
    x"e84088b8",
    x"54427fff",
    x"c45fffff",
    x"54217fff",
    x"c43ffffc",
    x"e3c00000",
    x"579c7ff4",
    x"2fdc0000",
    x"2e9c0004",
    x"2ebc0008",
    x"ee980000",
    x"eaa00001",
    x"2eb40000",
    x"00202a10",
    x"e7e0000a",
    x"e8200010",
    x"e7ffffef",
    x"56b50001",
    x"c01ffffa",
    x"0fdc0000",
    x"0e9c0004",
    x"0ebc0008",
    x"579c000c",
    x"e3c00000",
    x"579c7ffc",
    x"2fdc0000",
    x"e7e00004",
    x"0fdc0000",
    x"579c0004",
    x"e3c00000",
    x"579c7ffc",
    x"2e9c0000",
    x"0dbf00e8",
    x"0e3f00d4",
    x"0e5f00d4",
    x"00210068",
    x"00210272",
    x"ec478478",
    x"00410472",
    x"ec67f000",
    x"00420670",
    x"02830473",
    x"01ad2872",
    x"edc80002",
    x"41ce0000",
    x"ea000168",
    x"84700001",
    x"00630068",
    x"006d0672",
    x"0c5f00a0",
    x"00420671",
    x"e9e00280",
    x"846f0001",
    x"00630068",
    x"006d0672",
    x"0c3f0084",
    x"00210671",
    x"00600010",
    x"00800010",
    x"e9200000",
    x"00a30672",
    x"00c40872",
    x"55290001",
    x"00830872",
    x"00650c71",
    x"00a50c70",
    x"00840870",
    x"00630270",
    x"01492219",
    x"00840470",
    x"00a52464",
    x"cca00003",
    x"c95ffff4",
    x"e9200000",
    x"89290001",
    x"252e0000",
    x"55ce0001",
    x"55ef7fff",
    x"00211a70",
    x"ddffffea",
    x"56107fff",
    x"00421a70",
    x"de1fffe1",
    x"0e9c0000",
    x"579c0004",
    x"e3c00000",
    x"0000007f",
    x"40800000",
    x"bf9403b1",
    x"be8ef344",
    x"3be56042",
    x"000006b8",
    x"676f7270",
    x"006d6172",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000",
    x"00000000"
  );

  signal s_is_valid_wb_request : std_logic;
begin
  -- Wishbone control logic.
  s_is_valid_wb_request <= i_wb_cyc and i_wb_stb;

  -- We always ack and never stall - we're that fast ;-)
  process(i_clk)
  begin
    if rising_edge(i_clk) then
      o_wb_dat <= C_ROM_ARRAY(to_integer(unsigned(i_wb_adr(C_ADDR_BITS+1 downto 2))));
      o_wb_ack <= s_is_valid_wb_request;
    end if;
  end process;
  o_wb_stall <= '0';
end rtl;
