----------------------------------------------------------------------------------------------------
-- Copyright (c) 2019 Marcus Geelnard
--
-- This software is provided 'as-is', without any express or implied warranty. In no event will the
-- authors be held liable for any damages arising from the use of this software.
--
-- Permission is granted to anyone to use this software for any purpose, including commercial
-- applications, and to alter it and redistribute it freely, subject to the following restrictions:
--
--  1. The origin of this software must not be misrepresented; you must not claim that you wrote
--     the original software. If you use this software in a product, an acknowledgment in the
--     product documentation would be appreciated but is not required.
--
--  2. Altered source versions must be plainly marked as such, and must not be misrepresented as
--     being the original software.
--
--  3. This notice may not be removed or altered from any source distribution.
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
-- This is a single-ported ROM (Wishbone B4 pipelined interface).
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
  port(
    -- Control signals.
    i_clk : in std_logic;

    -- Wishbone memory interface (b4 pipelined slave).
    -- See: https://cdn.opencores.org/downloads/wbspec_b4.pdf
    i_wb_cyc : in std_logic;
    i_wb_stb : in std_logic;
    i_wb_adr : in std_logic_vector(31 downto 2);
    o_wb_dat : out std_logic_vector(31 downto 0);
    o_wb_ack : out std_logic;
    o_wb_stall : out std_logic
  );
end rom;

architecture rtl of rom is
  constant C_ADDR_BITS : positive := 10;

  signal s_is_valid_wb_request : std_logic;
  signal s_rom_addr : std_logic_vector(C_ADDR_BITS-1 downto 0);
begin
  -- Wishbone control logic.
  s_is_valid_wb_request <= i_wb_cyc and i_wb_stb;

  -- We always ack and never stall - we're that fast ;-)
  process(i_clk)
  begin
    if rising_edge(i_clk) then
      o_wb_ack <= s_is_valid_wb_request;
    end if;
  end process;
  o_wb_stall <= '0';

  -- Actual ROM.
  s_rom_addr <= i_wb_adr(C_ADDR_BITS+1 downto 2);

  process(i_clk)
  begin
    if rising_edge(i_clk) then
      case s_rom_addr is
        when 10x"0" => o_wb_dat <= x"00000000";
        when 10x"1" => o_wb_dat <= x"00000000";
        when 10x"2" => o_wb_dat <= x"00000000";
        when 10x"3" => o_wb_dat <= x"00000000";
        when 10x"4" => o_wb_dat <= x"00000000";
        when 10x"5" => o_wb_dat <= x"00000000";
        when 10x"6" => o_wb_dat <= x"00000000";
        when 10x"7" => o_wb_dat <= x"00000000";
        when 10x"8" => o_wb_dat <= x"00000000";
        when 10x"9" => o_wb_dat <= x"00000000";
        when 10x"a" => o_wb_dat <= x"00000000";
        when 10x"b" => o_wb_dat <= x"00000000";
        when 10x"c" => o_wb_dat <= x"00000000";
        when 10x"d" => o_wb_dat <= x"00000000";
        when 10x"e" => o_wb_dat <= x"00000000";
        when 10x"f" => o_wb_dat <= x"00000000";
        when 10x"10" => o_wb_dat <= x"00000000";
        when 10x"11" => o_wb_dat <= x"00000000";
        when 10x"12" => o_wb_dat <= x"00000000";
        when 10x"13" => o_wb_dat <= x"00000000";
        when 10x"14" => o_wb_dat <= x"00000000";
        when 10x"15" => o_wb_dat <= x"00000000";
        when 10x"16" => o_wb_dat <= x"00000000";
        when 10x"17" => o_wb_dat <= x"00000000";
        when 10x"18" => o_wb_dat <= x"00000000";
        when 10x"19" => o_wb_dat <= x"00000000";
        when 10x"1a" => o_wb_dat <= x"00000000";
        when 10x"1b" => o_wb_dat <= x"00000000";
        when 10x"1c" => o_wb_dat <= x"00000000";
        when 10x"1d" => o_wb_dat <= x"00000000";
        when 10x"1e" => o_wb_dat <= x"00000000";
        when 10x"1f" => o_wb_dat <= x"00000000";
        when 10x"20" => o_wb_dat <= x"00000000";
        when 10x"21" => o_wb_dat <= x"00000000";
        when 10x"22" => o_wb_dat <= x"00000000";
        when 10x"23" => o_wb_dat <= x"00000000";
        when 10x"24" => o_wb_dat <= x"00000000";
        when 10x"25" => o_wb_dat <= x"00000000";
        when 10x"26" => o_wb_dat <= x"00000000";
        when 10x"27" => o_wb_dat <= x"00000000";
        when 10x"28" => o_wb_dat <= x"00000000";
        when 10x"29" => o_wb_dat <= x"00000000";
        when 10x"2a" => o_wb_dat <= x"00000000";
        when 10x"2b" => o_wb_dat <= x"00000000";
        when 10x"2c" => o_wb_dat <= x"00000000";
        when 10x"2d" => o_wb_dat <= x"00000000";
        when 10x"2e" => o_wb_dat <= x"00000000";
        when 10x"2f" => o_wb_dat <= x"00000000";
        when 10x"30" => o_wb_dat <= x"00000000";
        when 10x"31" => o_wb_dat <= x"00000000";
        when 10x"32" => o_wb_dat <= x"00000000";
        when 10x"33" => o_wb_dat <= x"00000000";
        when 10x"34" => o_wb_dat <= x"00000000";
        when 10x"35" => o_wb_dat <= x"00000000";
        when 10x"36" => o_wb_dat <= x"00000000";
        when 10x"37" => o_wb_dat <= x"00000000";
        when 10x"38" => o_wb_dat <= x"00000000";
        when 10x"39" => o_wb_dat <= x"00000000";
        when 10x"3a" => o_wb_dat <= x"00000000";
        when 10x"3b" => o_wb_dat <= x"00000000";
        when 10x"3c" => o_wb_dat <= x"00000000";
        when 10x"3d" => o_wb_dat <= x"00000000";
        when 10x"3e" => o_wb_dat <= x"00000000";
        when 10x"3f" => o_wb_dat <= x"00000000";
        when 10x"40" => o_wb_dat <= x"00000000";
        when 10x"41" => o_wb_dat <= x"00000000";
        when 10x"42" => o_wb_dat <= x"00000000";
        when 10x"43" => o_wb_dat <= x"00000000";
        when 10x"44" => o_wb_dat <= x"00000000";
        when 10x"45" => o_wb_dat <= x"00000000";
        when 10x"46" => o_wb_dat <= x"00000000";
        when 10x"47" => o_wb_dat <= x"00000000";
        when 10x"48" => o_wb_dat <= x"00000000";
        when 10x"49" => o_wb_dat <= x"00000000";
        when 10x"4a" => o_wb_dat <= x"00000000";
        when 10x"4b" => o_wb_dat <= x"00000000";
        when 10x"4c" => o_wb_dat <= x"00000000";
        when 10x"4d" => o_wb_dat <= x"00000000";
        when 10x"4e" => o_wb_dat <= x"00000000";
        when 10x"4f" => o_wb_dat <= x"00000000";
        when 10x"50" => o_wb_dat <= x"00000000";
        when 10x"51" => o_wb_dat <= x"00000000";
        when 10x"52" => o_wb_dat <= x"00000000";
        when 10x"53" => o_wb_dat <= x"00000000";
        when 10x"54" => o_wb_dat <= x"00000000";
        when 10x"55" => o_wb_dat <= x"00000000";
        when 10x"56" => o_wb_dat <= x"00000000";
        when 10x"57" => o_wb_dat <= x"00000000";
        when 10x"58" => o_wb_dat <= x"00000000";
        when 10x"59" => o_wb_dat <= x"00000000";
        when 10x"5a" => o_wb_dat <= x"00000000";
        when 10x"5b" => o_wb_dat <= x"00000000";
        when 10x"5c" => o_wb_dat <= x"00000000";
        when 10x"5d" => o_wb_dat <= x"00000000";
        when 10x"5e" => o_wb_dat <= x"00000000";
        when 10x"5f" => o_wb_dat <= x"00000000";
        when 10x"60" => o_wb_dat <= x"00000000";
        when 10x"61" => o_wb_dat <= x"00000000";
        when 10x"62" => o_wb_dat <= x"00000000";
        when 10x"63" => o_wb_dat <= x"00000000";
        when 10x"64" => o_wb_dat <= x"00000000";
        when 10x"65" => o_wb_dat <= x"00000000";
        when 10x"66" => o_wb_dat <= x"00000000";
        when 10x"67" => o_wb_dat <= x"00000000";
        when 10x"68" => o_wb_dat <= x"00000000";
        when 10x"69" => o_wb_dat <= x"00000000";
        when 10x"6a" => o_wb_dat <= x"00000000";
        when 10x"6b" => o_wb_dat <= x"00000000";
        when 10x"6c" => o_wb_dat <= x"00000000";
        when 10x"6d" => o_wb_dat <= x"00000000";
        when 10x"6e" => o_wb_dat <= x"00000000";
        when 10x"6f" => o_wb_dat <= x"00000000";
        when 10x"70" => o_wb_dat <= x"00000000";
        when 10x"71" => o_wb_dat <= x"00000000";
        when 10x"72" => o_wb_dat <= x"00000000";
        when 10x"73" => o_wb_dat <= x"00000000";
        when 10x"74" => o_wb_dat <= x"00000000";
        when 10x"75" => o_wb_dat <= x"00000000";
        when 10x"76" => o_wb_dat <= x"00000000";
        when 10x"77" => o_wb_dat <= x"00000000";
        when 10x"78" => o_wb_dat <= x"00000000";
        when 10x"79" => o_wb_dat <= x"00000000";
        when 10x"7a" => o_wb_dat <= x"00000000";
        when 10x"7b" => o_wb_dat <= x"00000000";
        when 10x"7c" => o_wb_dat <= x"00000000";
        when 10x"7d" => o_wb_dat <= x"00000000";
        when 10x"7e" => o_wb_dat <= x"00000000";
        when 10x"7f" => o_wb_dat <= x"00000000";
        when 10x"80" => o_wb_dat <= x"579c7ffc";
        when 10x"81" => o_wb_dat <= x"2fdc0000";
        when 10x"82" => o_wb_dat <= x"e7e00005";
        when 10x"83" => o_wb_dat <= x"e7e0005e";
        when 10x"84" => o_wb_dat <= x"0fdc0000";
        when 10x"85" => o_wb_dat <= x"579c0004";
        when 10x"86" => o_wb_dat <= x"e3c00000";
        when 10x"87" => o_wb_dat <= x"579c7ffc";
        when 10x"88" => o_wb_dat <= x"2fbc0000";
        when 10x"89" => o_wb_dat <= x"ed680000";
        when 10x"8a" => o_wb_dat <= x"416b0000";
        when 10x"8b" => o_wb_dat <= x"ed90400a";
        when 10x"8c" => o_wb_dat <= x"418c0555";
        when 10x"8d" => o_wb_dat <= x"2d8b0000";
        when 10x"8e" => o_wb_dat <= x"ed90a000";
        when 10x"8f" => o_wb_dat <= x"418c0002";
        when 10x"90" => o_wb_dat <= x"2d8b0004";
        when 10x"91" => o_wb_dat <= x"ed90c000";
        when 10x"92" => o_wb_dat <= x"418c0001";
        when 10x"93" => o_wb_dat <= x"2d8b0008";
        when 10x"94" => o_wb_dat <= x"ed8c0000";
        when 10x"95" => o_wb_dat <= x"418c00ff";
        when 10x"96" => o_wb_dat <= x"2d8b000c";
        when 10x"97" => o_wb_dat <= x"556b0010";
        when 10x"98" => o_wb_dat <= x"e8200064";
        when 10x"99" => o_wb_dat <= x"e8400032";
        when 10x"9a" => o_wb_dat <= x"e8600000";
        when 10x"9b" => o_wb_dat <= x"e8800002";
        when 10x"9c" => o_wb_dat <= x"e8a00003";
        when 10x"9d" => o_wb_dat <= x"e8c00001";
        when 10x"9e" => o_wb_dat <= x"edffe000";
        when 10x"9f" => o_wb_dat <= x"2deb0000";
        when 10x"a0" => o_wb_dat <= x"e9c00001";
        when 10x"a1" => o_wb_dat <= x"88e30010";
        when 10x"a2" => o_wb_dat <= x"89020008";
        when 10x"a3" => o_wb_dat <= x"00e71010";
        when 10x"a4" => o_wb_dat <= x"00e70210";
        when 10x"a5" => o_wb_dat <= x"00e71e10";
        when 10x"a6" => o_wb_dat <= x"00eb1d0b";
        when 10x"a7" => o_wb_dat <= x"00210815";
        when 10x"a8" => o_wb_dat <= x"6ce100ff";
        when 10x"a9" => o_wb_dat <= x"0100021b";
        when 10x"aa" => o_wb_dat <= x"00e71012";
        when 10x"ab" => o_wb_dat <= x"c8e00003";
        when 10x"ac" => o_wb_dat <= x"00840016";
        when 10x"ad" => o_wb_dat <= x"00210815";
        when 10x"ae" => o_wb_dat <= x"00420a15";
        when 10x"af" => o_wb_dat <= x"6ce200ff";
        when 10x"b0" => o_wb_dat <= x"0100041b";
        when 10x"b1" => o_wb_dat <= x"00e71012";
        when 10x"b2" => o_wb_dat <= x"c8e00003";
        when 10x"b3" => o_wb_dat <= x"00a50016";
        when 10x"b4" => o_wb_dat <= x"00420a15";
        when 10x"b5" => o_wb_dat <= x"00630c15";
        when 10x"b6" => o_wb_dat <= x"6ce300ff";
        when 10x"b7" => o_wb_dat <= x"0100061b";
        when 10x"b8" => o_wb_dat <= x"00e71012";
        when 10x"b9" => o_wb_dat <= x"c8e00003";
        when 10x"ba" => o_wb_dat <= x"00c60016";
        when 10x"bb" => o_wb_dat <= x"00630c15";
        when 10x"bc" => o_wb_dat <= x"55ce0001";
        when 10x"bd" => o_wb_dat <= x"60ee0100";
        when 10x"be" => o_wb_dat <= x"c8ffffe3";
        when 10x"bf" => o_wb_dat <= x"556b0400";
        when 10x"c0" => o_wb_dat <= x"ec2a0000";
        when 10x"c1" => o_wb_dat <= x"ec500000";
        when 10x"c2" => o_wb_dat <= x"40420400";
        when 10x"c3" => o_wb_dat <= x"2c2b0000";
        when 10x"c4" => o_wb_dat <= x"2c4b0004";
        when 10x"c5" => o_wb_dat <= x"ed908000";
        when 10x"c6" => o_wb_dat <= x"418c0780";
        when 10x"c7" => o_wb_dat <= x"2d8b0008";
        when 10x"c8" => o_wb_dat <= x"556b000c";
        when 10x"c9" => o_wb_dat <= x"e3e00004";
        when 10x"ca" => o_wb_dat <= x"2c2b0000";
        when 10x"cb" => o_wb_dat <= x"2c4b0004";
        when 10x"cc" => o_wb_dat <= x"556b0008";
        when 10x"cd" => o_wb_dat <= x"54210003";
        when 10x"ce" => o_wb_dat <= x"544200a0";
        when 10x"cf" => o_wb_dat <= x"49a13fff";
        when 10x"d0" => o_wb_dat <= x"65ad0438";
        when 10x"d1" => o_wb_dat <= x"c9bffff9";
        when 10x"d2" => o_wb_dat <= x"ed8a000f";
        when 10x"d3" => o_wb_dat <= x"418c07ff";
        when 10x"d4" => o_wb_dat <= x"2d8b0000";
        when 10x"d5" => o_wb_dat <= x"ed280002";
        when 10x"d6" => o_wb_dat <= x"41290000";
        when 10x"d7" => o_wb_dat <= x"01400000";
        when 10x"d8" => o_wb_dat <= x"e960e100";
        when 10x"d9" => o_wb_dat <= x"03aa161d";
        when 10x"da" => o_wb_dat <= x"017d1616";
        when 10x"db" => o_wb_dat <= x"2c098004";
        when 10x"dc" => o_wb_dat <= x"01293b07";
        when 10x"dd" => o_wb_dat <= x"c57ffffc";
        when 10x"de" => o_wb_dat <= x"0fbc0000";
        when 10x"df" => o_wb_dat <= x"579c0004";
        when 10x"e0" => o_wb_dat <= x"e3c00000";
        when 10x"e1" => o_wb_dat <= x"579c7ff4";
        when 10x"e2" => o_wb_dat <= x"2fdc0000";
        when 10x"e3" => o_wb_dat <= x"2e9c0004";
        when 10x"e4" => o_wb_dat <= x"2ebc0008";
        when 10x"e5" => o_wb_dat <= x"ee980000";
        when 10x"e6" => o_wb_dat <= x"eaa00001";
        when 10x"e7" => o_wb_dat <= x"2eb40060";
        when 10x"e8" => o_wb_dat <= x"0c340020";
        when 10x"e9" => o_wb_dat <= x"e7e002d9";
        when 10x"ea" => o_wb_dat <= x"00202a10";
        when 10x"eb" => o_wb_dat <= x"e7e00008";
        when 10x"ec" => o_wb_dat <= x"56b50001";
        when 10x"ed" => o_wb_dat <= x"c01ffffa";
        when 10x"ee" => o_wb_dat <= x"0fdc0000";
        when 10x"ef" => o_wb_dat <= x"0e9c0004";
        when 10x"f0" => o_wb_dat <= x"0ebc0008";
        when 10x"f1" => o_wb_dat <= x"579c000c";
        when 10x"f2" => o_wb_dat <= x"e3c00000";
        when 10x"f3" => o_wb_dat <= x"579c7ffc";
        when 10x"f4" => o_wb_dat <= x"2fdc0000";
        when 10x"f5" => o_wb_dat <= x"ec580000";
        when 10x"f6" => o_wb_dat <= x"0c420028";
        when 10x"f7" => o_wb_dat <= x"48420001";
        when 10x"f8" => o_wb_dat <= x"c0400003";
        when 10x"f9" => o_wb_dat <= x"e7e00043";
        when 10x"fa" => o_wb_dat <= x"c0000002";
        when 10x"fb" => o_wb_dat <= x"e7e00004";
        when 10x"fc" => o_wb_dat <= x"0fdc0000";
        when 10x"fd" => o_wb_dat <= x"579c0004";
        when 10x"fe" => o_wb_dat <= x"e3c00000";
        when 10x"ff" => o_wb_dat <= x"579c7ffc";
        when 10x"100" => o_wb_dat <= x"2e9c0000";
        when 10x"101" => o_wb_dat <= x"0dbf00e8";
        when 10x"102" => o_wb_dat <= x"0e3f00d4";
        when 10x"103" => o_wb_dat <= x"0e5f00d4";
        when 10x"104" => o_wb_dat <= x"00210068";
        when 10x"105" => o_wb_dat <= x"00210272";
        when 10x"106" => o_wb_dat <= x"ec478478";
        when 10x"107" => o_wb_dat <= x"00410472";
        when 10x"108" => o_wb_dat <= x"ec67f000";
        when 10x"109" => o_wb_dat <= x"00420670";
        when 10x"10a" => o_wb_dat <= x"02830473";
        when 10x"10b" => o_wb_dat <= x"01ad2872";
        when 10x"10c" => o_wb_dat <= x"edc80002";
        when 10x"10d" => o_wb_dat <= x"41ce0000";
        when 10x"10e" => o_wb_dat <= x"ea000168";
        when 10x"10f" => o_wb_dat <= x"84700001";
        when 10x"110" => o_wb_dat <= x"00630068";
        when 10x"111" => o_wb_dat <= x"006d0672";
        when 10x"112" => o_wb_dat <= x"0c5f00a0";
        when 10x"113" => o_wb_dat <= x"00420671";
        when 10x"114" => o_wb_dat <= x"e9e00280";
        when 10x"115" => o_wb_dat <= x"846f0001";
        when 10x"116" => o_wb_dat <= x"00630068";
        when 10x"117" => o_wb_dat <= x"006d0672";
        when 10x"118" => o_wb_dat <= x"0c3f0084";
        when 10x"119" => o_wb_dat <= x"00210671";
        when 10x"11a" => o_wb_dat <= x"00600010";
        when 10x"11b" => o_wb_dat <= x"00800010";
        when 10x"11c" => o_wb_dat <= x"e9200000";
        when 10x"11d" => o_wb_dat <= x"00a30672";
        when 10x"11e" => o_wb_dat <= x"00c40872";
        when 10x"11f" => o_wb_dat <= x"55290001";
        when 10x"120" => o_wb_dat <= x"00830872";
        when 10x"121" => o_wb_dat <= x"00650c71";
        when 10x"122" => o_wb_dat <= x"00a50c70";
        when 10x"123" => o_wb_dat <= x"00840870";
        when 10x"124" => o_wb_dat <= x"00630270";
        when 10x"125" => o_wb_dat <= x"01492219";
        when 10x"126" => o_wb_dat <= x"00840470";
        when 10x"127" => o_wb_dat <= x"00a52464";
        when 10x"128" => o_wb_dat <= x"cca00003";
        when 10x"129" => o_wb_dat <= x"c95ffff4";
        when 10x"12a" => o_wb_dat <= x"e9200000";
        when 10x"12b" => o_wb_dat <= x"89290001";
        when 10x"12c" => o_wb_dat <= x"252e0000";
        when 10x"12d" => o_wb_dat <= x"55ce0001";
        when 10x"12e" => o_wb_dat <= x"55ef7fff";
        when 10x"12f" => o_wb_dat <= x"00211a70";
        when 10x"130" => o_wb_dat <= x"ddffffea";
        when 10x"131" => o_wb_dat <= x"56107fff";
        when 10x"132" => o_wb_dat <= x"00421a70";
        when 10x"133" => o_wb_dat <= x"de1fffe1";
        when 10x"134" => o_wb_dat <= x"0e9c0000";
        when 10x"135" => o_wb_dat <= x"579c0004";
        when 10x"136" => o_wb_dat <= x"e3c00000";
        when 10x"137" => o_wb_dat <= x"0000007f";
        when 10x"138" => o_wb_dat <= x"40800000";
        when 10x"139" => o_wb_dat <= x"bf9403b1";
        when 10x"13a" => o_wb_dat <= x"be8ef344";
        when 10x"13b" => o_wb_dat <= x"3be56042";
        when 10x"13c" => o_wb_dat <= x"579c7ff8";
        when 10x"13d" => o_wb_dat <= x"2e9c0000";
        when 10x"13e" => o_wb_dat <= x"2ebc0004";
        when 10x"13f" => o_wb_dat <= x"00210215";
        when 10x"140" => o_wb_dat <= x"01a00000";
        when 10x"141" => o_wb_dat <= x"03a01a10";
        when 10x"142" => o_wb_dat <= x"544d7fff";
        when 10x"143" => o_wb_dat <= x"1c82ffff";
        when 10x"144" => o_wb_dat <= x"56bf0074";
        when 10x"145" => o_wb_dat <= x"ecc80002";
        when 10x"146" => o_wb_dat <= x"40c60000";
        when 10x"147" => o_wb_dat <= x"e9000168";
        when 10x"148" => o_wb_dat <= x"55087fff";
        when 10x"149" => o_wb_dat <= x"01280215";
        when 10x"14a" => o_wb_dat <= x"e8e00140";
        when 10x"14b" => o_wb_dat <= x"03ad0e1d";
        when 10x"14c" => o_wb_dat <= x"00fd0e16";
        when 10x"14d" => o_wb_dat <= x"00e48e15";
        when 10x"14e" => o_wb_dat <= x"02870287";
        when 10x"14f" => o_wb_dat <= x"0124a815";
        when 10x"150" => o_wb_dat <= x"490983ff";
        when 10x"151" => o_wb_dat <= x"0115d082";
        when 10x"152" => o_wb_dat <= x"00e7d140";
        when 10x"153" => o_wb_dat <= x"00279315";
        when 10x"154" => o_wb_dat <= x"2c268002";
        when 10x"155" => o_wb_dat <= x"00c61a87";
        when 10x"156" => o_wb_dat <= x"dcfffff5";
        when 10x"157" => o_wb_dat <= x"dd1ffff1";
        when 10x"158" => o_wb_dat <= x"ed580000";
        when 10x"159" => o_wb_dat <= x"0d8a0020";
        when 10x"15a" => o_wb_dat <= x"0d6a0020";
        when 10x"15b" => o_wb_dat <= x"016b1818";
        when 10x"15c" => o_wb_dat <= x"cd7ffffe";
        when 10x"15d" => o_wb_dat <= x"0e9c0000";
        when 10x"15e" => o_wb_dat <= x"0ebc0004";
        when 10x"15f" => o_wb_dat <= x"579c0008";
        when 10x"160" => o_wb_dat <= x"e3c00000";
        when 10x"161" => o_wb_dat <= x"00c90000";
        when 10x"162" => o_wb_dat <= x"025b0192";
        when 10x"163" => o_wb_dat <= x"03ed0324";
        when 10x"164" => o_wb_dat <= x"057f04b6";
        when 10x"165" => o_wb_dat <= x"07110648";
        when 10x"166" => o_wb_dat <= x"08a207d9";
        when 10x"167" => o_wb_dat <= x"0a33096a";
        when 10x"168" => o_wb_dat <= x"0bc40afb";
        when 10x"169" => o_wb_dat <= x"0d540c8c";
        when 10x"16a" => o_wb_dat <= x"0ee30e1c";
        when 10x"16b" => o_wb_dat <= x"10720fab";
        when 10x"16c" => o_wb_dat <= x"1201113a";
        when 10x"16d" => o_wb_dat <= x"138f12c8";
        when 10x"16e" => o_wb_dat <= x"151c1455";
        when 10x"16f" => o_wb_dat <= x"16a815e2";
        when 10x"170" => o_wb_dat <= x"1833176e";
        when 10x"171" => o_wb_dat <= x"19be18f9";
        when 10x"172" => o_wb_dat <= x"1b471a82";
        when 10x"173" => o_wb_dat <= x"1ccf1c0b";
        when 10x"174" => o_wb_dat <= x"1e571d93";
        when 10x"175" => o_wb_dat <= x"1fdd1f1a";
        when 10x"176" => o_wb_dat <= x"2161209f";
        when 10x"177" => o_wb_dat <= x"22e52223";
        when 10x"178" => o_wb_dat <= x"246723a6";
        when 10x"179" => o_wb_dat <= x"25e82528";
        when 10x"17a" => o_wb_dat <= x"276726a8";
        when 10x"17b" => o_wb_dat <= x"28e52826";
        when 10x"17c" => o_wb_dat <= x"2a6129a3";
        when 10x"17d" => o_wb_dat <= x"2bdc2b1f";
        when 10x"17e" => o_wb_dat <= x"2d552c99";
        when 10x"17f" => o_wb_dat <= x"2ecc2e11";
        when 10x"180" => o_wb_dat <= x"30412f87";
        when 10x"181" => o_wb_dat <= x"31b530fb";
        when 10x"182" => o_wb_dat <= x"3326326e";
        when 10x"183" => o_wb_dat <= x"349633df";
        when 10x"184" => o_wb_dat <= x"3604354d";
        when 10x"185" => o_wb_dat <= x"376f36ba";
        when 10x"186" => o_wb_dat <= x"38d93824";
        when 10x"187" => o_wb_dat <= x"3a40398c";
        when 10x"188" => o_wb_dat <= x"3ba53af2";
        when 10x"189" => o_wb_dat <= x"3d073c56";
        when 10x"18a" => o_wb_dat <= x"3e683db8";
        when 10x"18b" => o_wb_dat <= x"3fc53f17";
        when 10x"18c" => o_wb_dat <= x"41214073";
        when 10x"18d" => o_wb_dat <= x"427a41ce";
        when 10x"18e" => o_wb_dat <= x"43d04325";
        when 10x"18f" => o_wb_dat <= x"4524447a";
        when 10x"190" => o_wb_dat <= x"467545cd";
        when 10x"191" => o_wb_dat <= x"47c3471c";
        when 10x"192" => o_wb_dat <= x"490f4869";
        when 10x"193" => o_wb_dat <= x"4a5849b4";
        when 10x"194" => o_wb_dat <= x"4b9d4afb";
        when 10x"195" => o_wb_dat <= x"4ce04c3f";
        when 10x"196" => o_wb_dat <= x"4e204d81";
        when 10x"197" => o_wb_dat <= x"4f5d4ebf";
        when 10x"198" => o_wb_dat <= x"50974ffb";
        when 10x"199" => o_wb_dat <= x"51ce5133";
        when 10x"19a" => o_wb_dat <= x"53025268";
        when 10x"19b" => o_wb_dat <= x"5432539b";
        when 10x"19c" => o_wb_dat <= x"556054c9";
        when 10x"19d" => o_wb_dat <= x"568a55f5";
        when 10x"19e" => o_wb_dat <= x"57b0571d";
        when 10x"19f" => o_wb_dat <= x"58d35842";
        when 10x"1a0" => o_wb_dat <= x"59f35964";
        when 10x"1a1" => o_wb_dat <= x"5b0f5a82";
        when 10x"1a2" => o_wb_dat <= x"5c285b9c";
        when 10x"1a3" => o_wb_dat <= x"5d3e5cb3";
        when 10x"1a4" => o_wb_dat <= x"5e4f5dc7";
        when 10x"1a5" => o_wb_dat <= x"5f5d5ed7";
        when 10x"1a6" => o_wb_dat <= x"60685fe3";
        when 10x"1a7" => o_wb_dat <= x"616e60eb";
        when 10x"1a8" => o_wb_dat <= x"627161f0";
        when 10x"1a9" => o_wb_dat <= x"637062f1";
        when 10x"1aa" => o_wb_dat <= x"646c63ee";
        when 10x"1ab" => o_wb_dat <= x"656364e8";
        when 10x"1ac" => o_wb_dat <= x"665665dd";
        when 10x"1ad" => o_wb_dat <= x"674666cf";
        when 10x"1ae" => o_wb_dat <= x"683267bc";
        when 10x"1af" => o_wb_dat <= x"691968a6";
        when 10x"1b0" => o_wb_dat <= x"69fd698b";
        when 10x"1b1" => o_wb_dat <= x"6adc6a6d";
        when 10x"1b2" => o_wb_dat <= x"6bb76b4a";
        when 10x"1b3" => o_wb_dat <= x"6c8e6c23";
        when 10x"1b4" => o_wb_dat <= x"6d616cf8";
        when 10x"1b5" => o_wb_dat <= x"6e306dc9";
        when 10x"1b6" => o_wb_dat <= x"6efb6e96";
        when 10x"1b7" => o_wb_dat <= x"6fc16f5e";
        when 10x"1b8" => o_wb_dat <= x"70837022";
        when 10x"1b9" => o_wb_dat <= x"714070e2";
        when 10x"1ba" => o_wb_dat <= x"71f9719d";
        when 10x"1bb" => o_wb_dat <= x"72ae7254";
        when 10x"1bc" => o_wb_dat <= x"735e7307";
        when 10x"1bd" => o_wb_dat <= x"740a73b5";
        when 10x"1be" => o_wb_dat <= x"74b2745f";
        when 10x"1bf" => o_wb_dat <= x"75557504";
        when 10x"1c0" => o_wb_dat <= x"75f375a5";
        when 10x"1c1" => o_wb_dat <= x"768d7641";
        when 10x"1c2" => o_wb_dat <= x"772276d8";
        when 10x"1c3" => o_wb_dat <= x"77b3776b";
        when 10x"1c4" => o_wb_dat <= x"783f77fa";
        when 10x"1c5" => o_wb_dat <= x"78c77884";
        when 10x"1c6" => o_wb_dat <= x"794a7909";
        when 10x"1c7" => o_wb_dat <= x"79c87989";
        when 10x"1c8" => o_wb_dat <= x"7a417a05";
        when 10x"1c9" => o_wb_dat <= x"7ab67a7c";
        when 10x"1ca" => o_wb_dat <= x"7b267aee";
        when 10x"1cb" => o_wb_dat <= x"7b917b5c";
        when 10x"1cc" => o_wb_dat <= x"7bf87bc5";
        when 10x"1cd" => o_wb_dat <= x"7c597c29";
        when 10x"1ce" => o_wb_dat <= x"7cb67c88";
        when 10x"1cf" => o_wb_dat <= x"7d0e7ce3";
        when 10x"1d0" => o_wb_dat <= x"7d627d39";
        when 10x"1d1" => o_wb_dat <= x"7db07d89";
        when 10x"1d2" => o_wb_dat <= x"7dfa7dd5";
        when 10x"1d3" => o_wb_dat <= x"7e3e7e1d";
        when 10x"1d4" => o_wb_dat <= x"7e7e7e5f";
        when 10x"1d5" => o_wb_dat <= x"7eb97e9c";
        when 10x"1d6" => o_wb_dat <= x"7eef7ed5";
        when 10x"1d7" => o_wb_dat <= x"7f217f09";
        when 10x"1d8" => o_wb_dat <= x"7f4d7f37";
        when 10x"1d9" => o_wb_dat <= x"7f747f61";
        when 10x"1da" => o_wb_dat <= x"7f977f86";
        when 10x"1db" => o_wb_dat <= x"7fb47fa6";
        when 10x"1dc" => o_wb_dat <= x"7fcd7fc1";
        when 10x"1dd" => o_wb_dat <= x"7fe17fd8";
        when 10x"1de" => o_wb_dat <= x"7ff07fe9";
        when 10x"1df" => o_wb_dat <= x"7ff97ff5";
        when 10x"1e0" => o_wb_dat <= x"7ffe7ffd";
        when 10x"1e1" => o_wb_dat <= x"7ffe7fff";
        when 10x"1e2" => o_wb_dat <= x"7ff97ffd";
        when 10x"1e3" => o_wb_dat <= x"7ff07ff5";
        when 10x"1e4" => o_wb_dat <= x"7fe17fe9";
        when 10x"1e5" => o_wb_dat <= x"7fcd7fd8";
        when 10x"1e6" => o_wb_dat <= x"7fb47fc1";
        when 10x"1e7" => o_wb_dat <= x"7f977fa6";
        when 10x"1e8" => o_wb_dat <= x"7f747f86";
        when 10x"1e9" => o_wb_dat <= x"7f4d7f61";
        when 10x"1ea" => o_wb_dat <= x"7f217f37";
        when 10x"1eb" => o_wb_dat <= x"7eef7f09";
        when 10x"1ec" => o_wb_dat <= x"7eb97ed5";
        when 10x"1ed" => o_wb_dat <= x"7e7e7e9c";
        when 10x"1ee" => o_wb_dat <= x"7e3e7e5f";
        when 10x"1ef" => o_wb_dat <= x"7dfa7e1d";
        when 10x"1f0" => o_wb_dat <= x"7db07dd5";
        when 10x"1f1" => o_wb_dat <= x"7d627d89";
        when 10x"1f2" => o_wb_dat <= x"7d0e7d39";
        when 10x"1f3" => o_wb_dat <= x"7cb67ce3";
        when 10x"1f4" => o_wb_dat <= x"7c597c88";
        when 10x"1f5" => o_wb_dat <= x"7bf87c29";
        when 10x"1f6" => o_wb_dat <= x"7b917bc5";
        when 10x"1f7" => o_wb_dat <= x"7b267b5c";
        when 10x"1f8" => o_wb_dat <= x"7ab67aee";
        when 10x"1f9" => o_wb_dat <= x"7a417a7c";
        when 10x"1fa" => o_wb_dat <= x"79c87a05";
        when 10x"1fb" => o_wb_dat <= x"794a7989";
        when 10x"1fc" => o_wb_dat <= x"78c77909";
        when 10x"1fd" => o_wb_dat <= x"783f7884";
        when 10x"1fe" => o_wb_dat <= x"77b377fa";
        when 10x"1ff" => o_wb_dat <= x"7722776b";
        when 10x"200" => o_wb_dat <= x"768d76d8";
        when 10x"201" => o_wb_dat <= x"75f37641";
        when 10x"202" => o_wb_dat <= x"755575a5";
        when 10x"203" => o_wb_dat <= x"74b27504";
        when 10x"204" => o_wb_dat <= x"740a745f";
        when 10x"205" => o_wb_dat <= x"735e73b5";
        when 10x"206" => o_wb_dat <= x"72ae7307";
        when 10x"207" => o_wb_dat <= x"71f97254";
        when 10x"208" => o_wb_dat <= x"7140719d";
        when 10x"209" => o_wb_dat <= x"708370e2";
        when 10x"20a" => o_wb_dat <= x"6fc17022";
        when 10x"20b" => o_wb_dat <= x"6efb6f5e";
        when 10x"20c" => o_wb_dat <= x"6e306e96";
        when 10x"20d" => o_wb_dat <= x"6d616dc9";
        when 10x"20e" => o_wb_dat <= x"6c8e6cf8";
        when 10x"20f" => o_wb_dat <= x"6bb76c23";
        when 10x"210" => o_wb_dat <= x"6adc6b4a";
        when 10x"211" => o_wb_dat <= x"69fd6a6d";
        when 10x"212" => o_wb_dat <= x"6919698b";
        when 10x"213" => o_wb_dat <= x"683268a6";
        when 10x"214" => o_wb_dat <= x"674667bc";
        when 10x"215" => o_wb_dat <= x"665666cf";
        when 10x"216" => o_wb_dat <= x"656365dd";
        when 10x"217" => o_wb_dat <= x"646c64e8";
        when 10x"218" => o_wb_dat <= x"637063ee";
        when 10x"219" => o_wb_dat <= x"627162f1";
        when 10x"21a" => o_wb_dat <= x"616e61f0";
        when 10x"21b" => o_wb_dat <= x"606860eb";
        when 10x"21c" => o_wb_dat <= x"5f5d5fe3";
        when 10x"21d" => o_wb_dat <= x"5e4f5ed7";
        when 10x"21e" => o_wb_dat <= x"5d3e5dc7";
        when 10x"21f" => o_wb_dat <= x"5c285cb3";
        when 10x"220" => o_wb_dat <= x"5b0f5b9c";
        when 10x"221" => o_wb_dat <= x"59f35a82";
        when 10x"222" => o_wb_dat <= x"58d35964";
        when 10x"223" => o_wb_dat <= x"57b05842";
        when 10x"224" => o_wb_dat <= x"568a571d";
        when 10x"225" => o_wb_dat <= x"556055f5";
        when 10x"226" => o_wb_dat <= x"543254c9";
        when 10x"227" => o_wb_dat <= x"5302539b";
        when 10x"228" => o_wb_dat <= x"51ce5268";
        when 10x"229" => o_wb_dat <= x"50975133";
        when 10x"22a" => o_wb_dat <= x"4f5d4ffb";
        when 10x"22b" => o_wb_dat <= x"4e204ebf";
        when 10x"22c" => o_wb_dat <= x"4ce04d81";
        when 10x"22d" => o_wb_dat <= x"4b9d4c3f";
        when 10x"22e" => o_wb_dat <= x"4a584afb";
        when 10x"22f" => o_wb_dat <= x"490f49b4";
        when 10x"230" => o_wb_dat <= x"47c34869";
        when 10x"231" => o_wb_dat <= x"4675471c";
        when 10x"232" => o_wb_dat <= x"452445cd";
        when 10x"233" => o_wb_dat <= x"43d0447a";
        when 10x"234" => o_wb_dat <= x"427a4325";
        when 10x"235" => o_wb_dat <= x"412141ce";
        when 10x"236" => o_wb_dat <= x"3fc54073";
        when 10x"237" => o_wb_dat <= x"3e683f17";
        when 10x"238" => o_wb_dat <= x"3d073db8";
        when 10x"239" => o_wb_dat <= x"3ba53c56";
        when 10x"23a" => o_wb_dat <= x"3a403af2";
        when 10x"23b" => o_wb_dat <= x"38d9398c";
        when 10x"23c" => o_wb_dat <= x"376f3824";
        when 10x"23d" => o_wb_dat <= x"360436ba";
        when 10x"23e" => o_wb_dat <= x"3496354d";
        when 10x"23f" => o_wb_dat <= x"332633df";
        when 10x"240" => o_wb_dat <= x"31b5326e";
        when 10x"241" => o_wb_dat <= x"304130fb";
        when 10x"242" => o_wb_dat <= x"2ecc2f87";
        when 10x"243" => o_wb_dat <= x"2d552e11";
        when 10x"244" => o_wb_dat <= x"2bdc2c99";
        when 10x"245" => o_wb_dat <= x"2a612b1f";
        when 10x"246" => o_wb_dat <= x"28e529a3";
        when 10x"247" => o_wb_dat <= x"27672826";
        when 10x"248" => o_wb_dat <= x"25e826a8";
        when 10x"249" => o_wb_dat <= x"24672528";
        when 10x"24a" => o_wb_dat <= x"22e523a6";
        when 10x"24b" => o_wb_dat <= x"21612223";
        when 10x"24c" => o_wb_dat <= x"1fdd209f";
        when 10x"24d" => o_wb_dat <= x"1e571f1a";
        when 10x"24e" => o_wb_dat <= x"1ccf1d93";
        when 10x"24f" => o_wb_dat <= x"1b471c0b";
        when 10x"250" => o_wb_dat <= x"19be1a82";
        when 10x"251" => o_wb_dat <= x"183318f9";
        when 10x"252" => o_wb_dat <= x"16a8176e";
        when 10x"253" => o_wb_dat <= x"151c15e2";
        when 10x"254" => o_wb_dat <= x"138f1455";
        when 10x"255" => o_wb_dat <= x"120112c8";
        when 10x"256" => o_wb_dat <= x"1072113a";
        when 10x"257" => o_wb_dat <= x"0ee30fab";
        when 10x"258" => o_wb_dat <= x"0d540e1c";
        when 10x"259" => o_wb_dat <= x"0bc40c8c";
        when 10x"25a" => o_wb_dat <= x"0a330afb";
        when 10x"25b" => o_wb_dat <= x"08a2096a";
        when 10x"25c" => o_wb_dat <= x"071107d9";
        when 10x"25d" => o_wb_dat <= x"057f0648";
        when 10x"25e" => o_wb_dat <= x"03ed04b6";
        when 10x"25f" => o_wb_dat <= x"025b0324";
        when 10x"260" => o_wb_dat <= x"00c90192";
        when 10x"261" => o_wb_dat <= x"ff370000";
        when 10x"262" => o_wb_dat <= x"fda5fe6e";
        when 10x"263" => o_wb_dat <= x"fc13fcdc";
        when 10x"264" => o_wb_dat <= x"fa81fb4a";
        when 10x"265" => o_wb_dat <= x"f8eff9b8";
        when 10x"266" => o_wb_dat <= x"f75ef827";
        when 10x"267" => o_wb_dat <= x"f5cdf696";
        when 10x"268" => o_wb_dat <= x"f43cf505";
        when 10x"269" => o_wb_dat <= x"f2acf374";
        when 10x"26a" => o_wb_dat <= x"f11df1e4";
        when 10x"26b" => o_wb_dat <= x"ef8ef055";
        when 10x"26c" => o_wb_dat <= x"edffeec6";
        when 10x"26d" => o_wb_dat <= x"ec71ed38";
        when 10x"26e" => o_wb_dat <= x"eae4ebab";
        when 10x"26f" => o_wb_dat <= x"e958ea1e";
        when 10x"270" => o_wb_dat <= x"e7cde892";
        when 10x"271" => o_wb_dat <= x"e642e707";
        when 10x"272" => o_wb_dat <= x"e4b9e57e";
        when 10x"273" => o_wb_dat <= x"e331e3f5";
        when 10x"274" => o_wb_dat <= x"e1a9e26d";
        when 10x"275" => o_wb_dat <= x"e023e0e6";
        when 10x"276" => o_wb_dat <= x"de9fdf61";
        when 10x"277" => o_wb_dat <= x"dd1bdddd";
        when 10x"278" => o_wb_dat <= x"db99dc5a";
        when 10x"279" => o_wb_dat <= x"da18dad8";
        when 10x"27a" => o_wb_dat <= x"d899d958";
        when 10x"27b" => o_wb_dat <= x"d71bd7da";
        when 10x"27c" => o_wb_dat <= x"d59fd65d";
        when 10x"27d" => o_wb_dat <= x"d424d4e1";
        when 10x"27e" => o_wb_dat <= x"d2abd367";
        when 10x"27f" => o_wb_dat <= x"d134d1ef";
        when 10x"280" => o_wb_dat <= x"cfbfd079";
        when 10x"281" => o_wb_dat <= x"ce4bcf05";
        when 10x"282" => o_wb_dat <= x"ccdacd92";
        when 10x"283" => o_wb_dat <= x"cb6acc21";
        when 10x"284" => o_wb_dat <= x"c9fccab3";
        when 10x"285" => o_wb_dat <= x"c891c946";
        when 10x"286" => o_wb_dat <= x"c727c7dc";
        when 10x"287" => o_wb_dat <= x"c5c0c674";
        when 10x"288" => o_wb_dat <= x"c45bc50e";
        when 10x"289" => o_wb_dat <= x"c2f9c3aa";
        when 10x"28a" => o_wb_dat <= x"c198c248";
        when 10x"28b" => o_wb_dat <= x"c03bc0e9";
        when 10x"28c" => o_wb_dat <= x"bedfbf8d";
        when 10x"28d" => o_wb_dat <= x"bd86be32";
        when 10x"28e" => o_wb_dat <= x"bc30bcdb";
        when 10x"28f" => o_wb_dat <= x"badcbb86";
        when 10x"290" => o_wb_dat <= x"b98bba33";
        when 10x"291" => o_wb_dat <= x"b83db8e4";
        when 10x"292" => o_wb_dat <= x"b6f1b797";
        when 10x"293" => o_wb_dat <= x"b5a8b64c";
        when 10x"294" => o_wb_dat <= x"b463b505";
        when 10x"295" => o_wb_dat <= x"b320b3c1";
        when 10x"296" => o_wb_dat <= x"b1e0b27f";
        when 10x"297" => o_wb_dat <= x"b0a3b141";
        when 10x"298" => o_wb_dat <= x"af69b005";
        when 10x"299" => o_wb_dat <= x"ae32aecd";
        when 10x"29a" => o_wb_dat <= x"acfead98";
        when 10x"29b" => o_wb_dat <= x"abceac65";
        when 10x"29c" => o_wb_dat <= x"aaa0ab37";
        when 10x"29d" => o_wb_dat <= x"a976aa0b";
        when 10x"29e" => o_wb_dat <= x"a850a8e3";
        when 10x"29f" => o_wb_dat <= x"a72da7be";
        when 10x"2a0" => o_wb_dat <= x"a60da69c";
        when 10x"2a1" => o_wb_dat <= x"a4f1a57e";
        when 10x"2a2" => o_wb_dat <= x"a3d8a464";
        when 10x"2a3" => o_wb_dat <= x"a2c2a34d";
        when 10x"2a4" => o_wb_dat <= x"a1b1a239";
        when 10x"2a5" => o_wb_dat <= x"a0a3a129";
        when 10x"2a6" => o_wb_dat <= x"9f98a01d";
        when 10x"2a7" => o_wb_dat <= x"9e929f15";
        when 10x"2a8" => o_wb_dat <= x"9d8f9e10";
        when 10x"2a9" => o_wb_dat <= x"9c909d0f";
        when 10x"2aa" => o_wb_dat <= x"9b949c12";
        when 10x"2ab" => o_wb_dat <= x"9a9d9b18";
        when 10x"2ac" => o_wb_dat <= x"99aa9a23";
        when 10x"2ad" => o_wb_dat <= x"98ba9931";
        when 10x"2ae" => o_wb_dat <= x"97ce9844";
        when 10x"2af" => o_wb_dat <= x"96e7975a";
        when 10x"2b0" => o_wb_dat <= x"96039675";
        when 10x"2b1" => o_wb_dat <= x"95249593";
        when 10x"2b2" => o_wb_dat <= x"944994b6";
        when 10x"2b3" => o_wb_dat <= x"937293dd";
        when 10x"2b4" => o_wb_dat <= x"929f9308";
        when 10x"2b5" => o_wb_dat <= x"91d09237";
        when 10x"2b6" => o_wb_dat <= x"9105916a";
        when 10x"2b7" => o_wb_dat <= x"903f90a2";
        when 10x"2b8" => o_wb_dat <= x"8f7d8fde";
        when 10x"2b9" => o_wb_dat <= x"8ec08f1e";
        when 10x"2ba" => o_wb_dat <= x"8e078e63";
        when 10x"2bb" => o_wb_dat <= x"8d528dac";
        when 10x"2bc" => o_wb_dat <= x"8ca28cf9";
        when 10x"2bd" => o_wb_dat <= x"8bf68c4b";
        when 10x"2be" => o_wb_dat <= x"8b4e8ba1";
        when 10x"2bf" => o_wb_dat <= x"8aab8afc";
        when 10x"2c0" => o_wb_dat <= x"8a0d8a5b";
        when 10x"2c1" => o_wb_dat <= x"897389bf";
        when 10x"2c2" => o_wb_dat <= x"88de8928";
        when 10x"2c3" => o_wb_dat <= x"884d8895";
        when 10x"2c4" => o_wb_dat <= x"87c18806";
        when 10x"2c5" => o_wb_dat <= x"8739877c";
        when 10x"2c6" => o_wb_dat <= x"86b686f7";
        when 10x"2c7" => o_wb_dat <= x"86388677";
        when 10x"2c8" => o_wb_dat <= x"85bf85fb";
        when 10x"2c9" => o_wb_dat <= x"854a8584";
        when 10x"2ca" => o_wb_dat <= x"84da8512";
        when 10x"2cb" => o_wb_dat <= x"846f84a4";
        when 10x"2cc" => o_wb_dat <= x"8408843b";
        when 10x"2cd" => o_wb_dat <= x"83a783d7";
        when 10x"2ce" => o_wb_dat <= x"834a8378";
        when 10x"2cf" => o_wb_dat <= x"82f2831d";
        when 10x"2d0" => o_wb_dat <= x"829e82c7";
        when 10x"2d1" => o_wb_dat <= x"82508277";
        when 10x"2d2" => o_wb_dat <= x"8206822b";
        when 10x"2d3" => o_wb_dat <= x"81c281e3";
        when 10x"2d4" => o_wb_dat <= x"818281a1";
        when 10x"2d5" => o_wb_dat <= x"81478164";
        when 10x"2d6" => o_wb_dat <= x"8111812b";
        when 10x"2d7" => o_wb_dat <= x"80df80f7";
        when 10x"2d8" => o_wb_dat <= x"80b380c9";
        when 10x"2d9" => o_wb_dat <= x"808c809f";
        when 10x"2da" => o_wb_dat <= x"8069807a";
        when 10x"2db" => o_wb_dat <= x"804c805a";
        when 10x"2dc" => o_wb_dat <= x"8033803f";
        when 10x"2dd" => o_wb_dat <= x"801f8028";
        when 10x"2de" => o_wb_dat <= x"80108017";
        when 10x"2df" => o_wb_dat <= x"8007800b";
        when 10x"2e0" => o_wb_dat <= x"80028003";
        when 10x"2e1" => o_wb_dat <= x"80028001";
        when 10x"2e2" => o_wb_dat <= x"80078003";
        when 10x"2e3" => o_wb_dat <= x"8010800b";
        when 10x"2e4" => o_wb_dat <= x"801f8017";
        when 10x"2e5" => o_wb_dat <= x"80338028";
        when 10x"2e6" => o_wb_dat <= x"804c803f";
        when 10x"2e7" => o_wb_dat <= x"8069805a";
        when 10x"2e8" => o_wb_dat <= x"808c807a";
        when 10x"2e9" => o_wb_dat <= x"80b3809f";
        when 10x"2ea" => o_wb_dat <= x"80df80c9";
        when 10x"2eb" => o_wb_dat <= x"811180f7";
        when 10x"2ec" => o_wb_dat <= x"8147812b";
        when 10x"2ed" => o_wb_dat <= x"81828164";
        when 10x"2ee" => o_wb_dat <= x"81c281a1";
        when 10x"2ef" => o_wb_dat <= x"820681e3";
        when 10x"2f0" => o_wb_dat <= x"8250822b";
        when 10x"2f1" => o_wb_dat <= x"829e8277";
        when 10x"2f2" => o_wb_dat <= x"82f282c7";
        when 10x"2f3" => o_wb_dat <= x"834a831d";
        when 10x"2f4" => o_wb_dat <= x"83a78378";
        when 10x"2f5" => o_wb_dat <= x"840883d7";
        when 10x"2f6" => o_wb_dat <= x"846f843b";
        when 10x"2f7" => o_wb_dat <= x"84da84a4";
        when 10x"2f8" => o_wb_dat <= x"854a8512";
        when 10x"2f9" => o_wb_dat <= x"85bf8584";
        when 10x"2fa" => o_wb_dat <= x"863885fb";
        when 10x"2fb" => o_wb_dat <= x"86b68677";
        when 10x"2fc" => o_wb_dat <= x"873986f7";
        when 10x"2fd" => o_wb_dat <= x"87c1877c";
        when 10x"2fe" => o_wb_dat <= x"884d8806";
        when 10x"2ff" => o_wb_dat <= x"88de8895";
        when 10x"300" => o_wb_dat <= x"89738928";
        when 10x"301" => o_wb_dat <= x"8a0d89bf";
        when 10x"302" => o_wb_dat <= x"8aab8a5b";
        when 10x"303" => o_wb_dat <= x"8b4e8afc";
        when 10x"304" => o_wb_dat <= x"8bf68ba1";
        when 10x"305" => o_wb_dat <= x"8ca28c4b";
        when 10x"306" => o_wb_dat <= x"8d528cf9";
        when 10x"307" => o_wb_dat <= x"8e078dac";
        when 10x"308" => o_wb_dat <= x"8ec08e63";
        when 10x"309" => o_wb_dat <= x"8f7d8f1e";
        when 10x"30a" => o_wb_dat <= x"903f8fde";
        when 10x"30b" => o_wb_dat <= x"910590a2";
        when 10x"30c" => o_wb_dat <= x"91d0916a";
        when 10x"30d" => o_wb_dat <= x"929f9237";
        when 10x"30e" => o_wb_dat <= x"93729308";
        when 10x"30f" => o_wb_dat <= x"944993dd";
        when 10x"310" => o_wb_dat <= x"952494b6";
        when 10x"311" => o_wb_dat <= x"96039593";
        when 10x"312" => o_wb_dat <= x"96e79675";
        when 10x"313" => o_wb_dat <= x"97ce975a";
        when 10x"314" => o_wb_dat <= x"98ba9844";
        when 10x"315" => o_wb_dat <= x"99aa9931";
        when 10x"316" => o_wb_dat <= x"9a9d9a23";
        when 10x"317" => o_wb_dat <= x"9b949b18";
        when 10x"318" => o_wb_dat <= x"9c909c12";
        when 10x"319" => o_wb_dat <= x"9d8f9d0f";
        when 10x"31a" => o_wb_dat <= x"9e929e10";
        when 10x"31b" => o_wb_dat <= x"9f989f15";
        when 10x"31c" => o_wb_dat <= x"a0a3a01d";
        when 10x"31d" => o_wb_dat <= x"a1b1a129";
        when 10x"31e" => o_wb_dat <= x"a2c2a239";
        when 10x"31f" => o_wb_dat <= x"a3d8a34d";
        when 10x"320" => o_wb_dat <= x"a4f1a464";
        when 10x"321" => o_wb_dat <= x"a60da57e";
        when 10x"322" => o_wb_dat <= x"a72da69c";
        when 10x"323" => o_wb_dat <= x"a850a7be";
        when 10x"324" => o_wb_dat <= x"a976a8e3";
        when 10x"325" => o_wb_dat <= x"aaa0aa0b";
        when 10x"326" => o_wb_dat <= x"abceab37";
        when 10x"327" => o_wb_dat <= x"acfeac65";
        when 10x"328" => o_wb_dat <= x"ae32ad98";
        when 10x"329" => o_wb_dat <= x"af69aecd";
        when 10x"32a" => o_wb_dat <= x"b0a3b005";
        when 10x"32b" => o_wb_dat <= x"b1e0b141";
        when 10x"32c" => o_wb_dat <= x"b320b27f";
        when 10x"32d" => o_wb_dat <= x"b463b3c1";
        when 10x"32e" => o_wb_dat <= x"b5a8b505";
        when 10x"32f" => o_wb_dat <= x"b6f1b64c";
        when 10x"330" => o_wb_dat <= x"b83db797";
        when 10x"331" => o_wb_dat <= x"b98bb8e4";
        when 10x"332" => o_wb_dat <= x"badcba33";
        when 10x"333" => o_wb_dat <= x"bc30bb86";
        when 10x"334" => o_wb_dat <= x"bd86bcdb";
        when 10x"335" => o_wb_dat <= x"bedfbe32";
        when 10x"336" => o_wb_dat <= x"c03bbf8d";
        when 10x"337" => o_wb_dat <= x"c198c0e9";
        when 10x"338" => o_wb_dat <= x"c2f9c248";
        when 10x"339" => o_wb_dat <= x"c45bc3aa";
        when 10x"33a" => o_wb_dat <= x"c5c0c50e";
        when 10x"33b" => o_wb_dat <= x"c727c674";
        when 10x"33c" => o_wb_dat <= x"c891c7dc";
        when 10x"33d" => o_wb_dat <= x"c9fcc946";
        when 10x"33e" => o_wb_dat <= x"cb6acab3";
        when 10x"33f" => o_wb_dat <= x"ccdacc21";
        when 10x"340" => o_wb_dat <= x"ce4bcd92";
        when 10x"341" => o_wb_dat <= x"cfbfcf05";
        when 10x"342" => o_wb_dat <= x"d134d079";
        when 10x"343" => o_wb_dat <= x"d2abd1ef";
        when 10x"344" => o_wb_dat <= x"d424d367";
        when 10x"345" => o_wb_dat <= x"d59fd4e1";
        when 10x"346" => o_wb_dat <= x"d71bd65d";
        when 10x"347" => o_wb_dat <= x"d899d7da";
        when 10x"348" => o_wb_dat <= x"da18d958";
        when 10x"349" => o_wb_dat <= x"db99dad8";
        when 10x"34a" => o_wb_dat <= x"dd1bdc5a";
        when 10x"34b" => o_wb_dat <= x"de9fdddd";
        when 10x"34c" => o_wb_dat <= x"e023df61";
        when 10x"34d" => o_wb_dat <= x"e1a9e0e6";
        when 10x"34e" => o_wb_dat <= x"e331e26d";
        when 10x"34f" => o_wb_dat <= x"e4b9e3f5";
        when 10x"350" => o_wb_dat <= x"e642e57e";
        when 10x"351" => o_wb_dat <= x"e7cde707";
        when 10x"352" => o_wb_dat <= x"e958e892";
        when 10x"353" => o_wb_dat <= x"eae4ea1e";
        when 10x"354" => o_wb_dat <= x"ec71ebab";
        when 10x"355" => o_wb_dat <= x"edffed38";
        when 10x"356" => o_wb_dat <= x"ef8eeec6";
        when 10x"357" => o_wb_dat <= x"f11df055";
        when 10x"358" => o_wb_dat <= x"f2acf1e4";
        when 10x"359" => o_wb_dat <= x"f43cf374";
        when 10x"35a" => o_wb_dat <= x"f5cdf505";
        when 10x"35b" => o_wb_dat <= x"f75ef696";
        when 10x"35c" => o_wb_dat <= x"f8eff827";
        when 10x"35d" => o_wb_dat <= x"fa81f9b8";
        when 10x"35e" => o_wb_dat <= x"fc13fb4a";
        when 10x"35f" => o_wb_dat <= x"fda5fcdc";
        when 10x"360" => o_wb_dat <= x"ff37fe6e";
        when 10x"361" => o_wb_dat <= x"e8200000";
        when 10x"362" => o_wb_dat <= x"e8400000";
        when 10x"363" => o_wb_dat <= x"e8600000";
        when 10x"364" => o_wb_dat <= x"e8800000";
        when 10x"365" => o_wb_dat <= x"e8a00000";
        when 10x"366" => o_wb_dat <= x"e8c00000";
        when 10x"367" => o_wb_dat <= x"e8e00000";
        when 10x"368" => o_wb_dat <= x"e9000000";
        when 10x"369" => o_wb_dat <= x"e9200000";
        when 10x"36a" => o_wb_dat <= x"e9400000";
        when 10x"36b" => o_wb_dat <= x"e9600000";
        when 10x"36c" => o_wb_dat <= x"e9800000";
        when 10x"36d" => o_wb_dat <= x"e9a00000";
        when 10x"36e" => o_wb_dat <= x"e9c00000";
        when 10x"36f" => o_wb_dat <= x"e9e00000";
        when 10x"370" => o_wb_dat <= x"ea000000";
        when 10x"371" => o_wb_dat <= x"ea200000";
        when 10x"372" => o_wb_dat <= x"ea400000";
        when 10x"373" => o_wb_dat <= x"ea600000";
        when 10x"374" => o_wb_dat <= x"ea800000";
        when 10x"375" => o_wb_dat <= x"eaa00000";
        when 10x"376" => o_wb_dat <= x"eac00000";
        when 10x"377" => o_wb_dat <= x"eae00000";
        when 10x"378" => o_wb_dat <= x"eb000000";
        when 10x"379" => o_wb_dat <= x"eb200000";
        when 10x"37a" => o_wb_dat <= x"eb400000";
        when 10x"37b" => o_wb_dat <= x"eb600000";
        when 10x"37c" => o_wb_dat <= x"eb800000";
        when 10x"37d" => o_wb_dat <= x"eba00000";
        when 10x"37e" => o_wb_dat <= x"ebc00000";
        when 10x"37f" => o_wb_dat <= x"03a00000";
        when 10x"380" => o_wb_dat <= x"40208000";
        when 10x"381" => o_wb_dat <= x"40408000";
        when 10x"382" => o_wb_dat <= x"40608000";
        when 10x"383" => o_wb_dat <= x"40808000";
        when 10x"384" => o_wb_dat <= x"40a08000";
        when 10x"385" => o_wb_dat <= x"40c08000";
        when 10x"386" => o_wb_dat <= x"40e08000";
        when 10x"387" => o_wb_dat <= x"41008000";
        when 10x"388" => o_wb_dat <= x"41208000";
        when 10x"389" => o_wb_dat <= x"41408000";
        when 10x"38a" => o_wb_dat <= x"41608000";
        when 10x"38b" => o_wb_dat <= x"41808000";
        when 10x"38c" => o_wb_dat <= x"41a08000";
        when 10x"38d" => o_wb_dat <= x"41c08000";
        when 10x"38e" => o_wb_dat <= x"41e08000";
        when 10x"38f" => o_wb_dat <= x"42008000";
        when 10x"390" => o_wb_dat <= x"42208000";
        when 10x"391" => o_wb_dat <= x"42408000";
        when 10x"392" => o_wb_dat <= x"42608000";
        when 10x"393" => o_wb_dat <= x"42808000";
        when 10x"394" => o_wb_dat <= x"42a08000";
        when 10x"395" => o_wb_dat <= x"42c08000";
        when 10x"396" => o_wb_dat <= x"42e08000";
        when 10x"397" => o_wb_dat <= x"43008000";
        when 10x"398" => o_wb_dat <= x"43208000";
        when 10x"399" => o_wb_dat <= x"43408000";
        when 10x"39a" => o_wb_dat <= x"43608000";
        when 10x"39b" => o_wb_dat <= x"43808000";
        when 10x"39c" => o_wb_dat <= x"43a08000";
        when 10x"39d" => o_wb_dat <= x"43c08000";
        when 10x"39e" => o_wb_dat <= x"43e08000";
        when 10x"39f" => o_wb_dat <= x"ec380000";
        when 10x"3a0" => o_wb_dat <= x"0c21000c";
        when 10x"3a1" => o_wb_dat <= x"ef880000";
        when 10x"3a2" => o_wb_dat <= x"039c0215";
        when 10x"3a3" => o_wb_dat <= x"e8200001";
        when 10x"3a4" => o_wb_dat <= x"ec400001";
        when 10x"3a5" => o_wb_dat <= x"54420758";
        when 10x"3a6" => o_wb_dat <= x"ede00000";
        when 10x"3a7" => o_wb_dat <= x"e5e00080";
        when 10x"3a8" => o_wb_dat <= x"00000000";
        when 10x"3a9" => o_wb_dat <= x"00000000";
        when 10x"3aa" => o_wb_dat <= x"00000000";
        when 10x"3ab" => o_wb_dat <= x"00000000";
        when 10x"3ac" => o_wb_dat <= x"00000000";
        when 10x"3ad" => o_wb_dat <= x"e3e00000";
        when 10x"3ae" => o_wb_dat <= x"00000000";
        when 10x"3af" => o_wb_dat <= x"00000000";
        when 10x"3b0" => o_wb_dat <= x"00000000";
        when 10x"3b1" => o_wb_dat <= x"00000000";
        when 10x"3b2" => o_wb_dat <= x"00000000";
        when 10x"3b3" => o_wb_dat <= x"1c5f007c";
        when 10x"3b4" => o_wb_dat <= x"ec780000";
        when 10x"3b5" => o_wb_dat <= x"1c630040";
        when 10x"3b6" => o_wb_dat <= x"e8a00008";
        when 10x"3b7" => o_wb_dat <= x"4881000f";
        when 10x"3b8" => o_wb_dat <= x"8c210004";
        when 10x"3b9" => o_wb_dat <= x"00820805";
        when 10x"3ba" => o_wb_dat <= x"2c830000";
        when 10x"3bb" => o_wb_dat <= x"54630004";
        when 10x"3bc" => o_wb_dat <= x"54a57fff";
        when 10x"3bd" => o_wb_dat <= x"c0a00004";
        when 10x"3be" => o_wb_dat <= x"c43ffff9";
        when 10x"3bf" => o_wb_dat <= x"e8800000";
        when 10x"3c0" => o_wb_dat <= x"c03ffffa";
        when 10x"3c1" => o_wb_dat <= x"e3c00000";
        when 10x"3c2" => o_wb_dat <= x"1c5f0040";
        when 10x"3c3" => o_wb_dat <= x"ec780000";
        when 10x"3c4" => o_wb_dat <= x"1c630040";
        when 10x"3c5" => o_wb_dat <= x"e8c0000a";
        when 10x"3c6" => o_wb_dat <= x"e8a00008";
        when 10x"3c7" => o_wb_dat <= x"00810c47";
        when 10x"3c8" => o_wb_dat <= x"00210c45";
        when 10x"3c9" => o_wb_dat <= x"00820805";
        when 10x"3ca" => o_wb_dat <= x"2c830000";
        when 10x"3cb" => o_wb_dat <= x"54630004";
        when 10x"3cc" => o_wb_dat <= x"54a57fff";
        when 10x"3cd" => o_wb_dat <= x"c0a00004";
        when 10x"3ce" => o_wb_dat <= x"c43ffff9";
        when 10x"3cf" => o_wb_dat <= x"e8800000";
        when 10x"3d0" => o_wb_dat <= x"c03ffffa";
        when 10x"3d1" => o_wb_dat <= x"e3c00000";
        when 10x"3d2" => o_wb_dat <= x"4f5b063f";
        when 10x"3d3" => o_wb_dat <= x"077d6d66";
        when 10x"3d4" => o_wb_dat <= x"7c776f7f";
        when 10x"3d5" => o_wb_dat <= x"71795e39";
        when 10x"3d6" => o_wb_dat <= x"00000f5c";
        when 10x"3d7" => o_wb_dat <= x"676f7270";
        when 10x"3d8" => o_wb_dat <= x"006d6172";
        when 10x"3d9" => o_wb_dat <= x"00000000";
        when 10x"3da" => o_wb_dat <= x"00000000";
        when 10x"3db" => o_wb_dat <= x"00000000";
        when 10x"3dc" => o_wb_dat <= x"00000000";
        when 10x"3dd" => o_wb_dat <= x"00000000";
        when 10x"3de" => o_wb_dat <= x"00000000";
        when 10x"3df" => o_wb_dat <= x"00000000";
        when 10x"3e0" => o_wb_dat <= x"00000000";
        when 10x"3e1" => o_wb_dat <= x"00000000";
        when 10x"3e2" => o_wb_dat <= x"00000000";
        when 10x"3e3" => o_wb_dat <= x"00000000";
        when 10x"3e4" => o_wb_dat <= x"00000000";
        when 10x"3e5" => o_wb_dat <= x"00000000";
        when 10x"3e6" => o_wb_dat <= x"00000000";
        when 10x"3e7" => o_wb_dat <= x"00000000";
        when 10x"3e8" => o_wb_dat <= x"00000000";
        when 10x"3e9" => o_wb_dat <= x"00000000";
        when 10x"3ea" => o_wb_dat <= x"00000000";
        when 10x"3eb" => o_wb_dat <= x"00000000";
        when 10x"3ec" => o_wb_dat <= x"00000000";
        when 10x"3ed" => o_wb_dat <= x"00000000";
        when 10x"3ee" => o_wb_dat <= x"00000000";
        when 10x"3ef" => o_wb_dat <= x"00000000";
        when 10x"3f0" => o_wb_dat <= x"00000000";
        when 10x"3f1" => o_wb_dat <= x"00000000";
        when 10x"3f2" => o_wb_dat <= x"00000000";
        when 10x"3f3" => o_wb_dat <= x"00000000";
        when 10x"3f4" => o_wb_dat <= x"00000000";
        when 10x"3f5" => o_wb_dat <= x"00000000";
        when 10x"3f6" => o_wb_dat <= x"00000000";
        when 10x"3f7" => o_wb_dat <= x"00000000";
        when 10x"3f8" => o_wb_dat <= x"00000000";
        when 10x"3f9" => o_wb_dat <= x"00000000";
        when 10x"3fa" => o_wb_dat <= x"00000000";
        when 10x"3fb" => o_wb_dat <= x"00000000";
        when 10x"3fc" => o_wb_dat <= x"00000000";
        when 10x"3fd" => o_wb_dat <= x"00000000";
        when 10x"3fe" => o_wb_dat <= x"00000000";
        when 10x"3ff" => o_wb_dat <= x"00000000";

        when others => o_wb_dat <= (others => '0');
      end case;
    end if;
  end process;
end rtl;
